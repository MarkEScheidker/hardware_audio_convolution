// Computer_System.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module Computer_System (
		input  wire        audio_ADCDAT,               //                audio.ADCDAT
		input  wire        audio_ADCLRCK,              //                     .ADCLRCK
		input  wire        audio_BCLK,                 //                     .BCLK
		output wire        audio_DACDAT,               //                     .DACDAT
		input  wire        audio_DACLRCK,              //                     .DACLRCK
		output wire        audio_pll_clk_clk,          //        audio_pll_clk.clk
		input  wire        audio_pll_ref_clk_clk,      //    audio_pll_ref_clk.clk
		input  wire        audio_pll_ref_reset_reset,  //  audio_pll_ref_reset.reset
		inout  wire        av_config_SDAT,             //            av_config.SDAT
		output wire        av_config_SCLK,             //                     .SCLK
		inout  wire [7:0]  char_lcd_DATA,              //             char_lcd.DATA
		output wire        char_lcd_ON,                //                     .ON
		output wire        char_lcd_BLON,              //                     .BLON
		output wire        char_lcd_EN,                //                     .EN
		output wire        char_lcd_RS,                //                     .RS
		output wire        char_lcd_RW,                //                     .RW
		inout  wire [31:0] expansion_jp5_export,       //        expansion_jp5.export
		output wire [22:0] flash_ADDR,                 //                flash.ADDR
		output wire        flash_CE_N,                 //                     .CE_N
		output wire        flash_OE_N,                 //                     .OE_N
		output wire        flash_WE_N,                 //                     .WE_N
		output wire        flash_RST_N,                //                     .RST_N
		inout  wire [7:0]  flash_DQ,                   //                     .DQ
		output wire [8:0]  green_leds_export,          //           green_leds.export
		output wire [31:0] hex3_hex0_export,           //            hex3_hex0.export
		output wire [31:0] hex7_hex4_export,           //            hex7_hex4.export
		output wire        irda_TXD,                   //                 irda.TXD
		input  wire        irda_RXD,                   //                     .RXD
		inout  wire        ps2_port_CLK,               //             ps2_port.CLK
		inout  wire        ps2_port_DAT,               //                     .DAT
		inout  wire        ps2_port_dual_CLK,          //        ps2_port_dual.CLK
		inout  wire        ps2_port_dual_DAT,          //                     .DAT
		input  wire [3:0]  pushbuttons_export,         //          pushbuttons.export
		output wire [17:0] red_leds_export,            //             red_leds.export
		inout  wire        sd_card_b_SD_cmd,           //              sd_card.b_SD_cmd
		inout  wire        sd_card_b_SD_dat,           //                     .b_SD_dat
		inout  wire        sd_card_b_SD_dat3,          //                     .b_SD_dat3
		output wire        sd_card_o_SD_clock,         //                     .o_SD_clock
		output wire [12:0] sdram_addr,                 //                sdram.addr
		output wire [1:0]  sdram_ba,                   //                     .ba
		output wire        sdram_cas_n,                //                     .cas_n
		output wire        sdram_cke,                  //                     .cke
		output wire        sdram_cs_n,                 //                     .cs_n
		inout  wire [31:0] sdram_dq,                   //                     .dq
		output wire [3:0]  sdram_dqm,                  //                     .dqm
		output wire        sdram_ras_n,                //                     .ras_n
		output wire        sdram_we_n,                 //                     .we_n
		output wire        sdram_clk_clk,              //            sdram_clk.clk
		input  wire        serial_port_RXD,            //          serial_port.RXD
		output wire        serial_port_TXD,            //                     .TXD
		input  wire [17:0] slider_switches_export,     //      slider_switches.export
		inout  wire [15:0] sram_DQ,                    //                 sram.DQ
		output wire [19:0] sram_ADDR,                  //                     .ADDR
		output wire        sram_LB_N,                  //                     .LB_N
		output wire        sram_UB_N,                  //                     .UB_N
		output wire        sram_CE_N,                  //                     .CE_N
		output wire        sram_OE_N,                  //                     .OE_N
		output wire        sram_WE_N,                  //                     .WE_N
		input  wire        system_pll_ref_clk_clk,     //   system_pll_ref_clk.clk
		input  wire        system_pll_ref_reset_reset, // system_pll_ref_reset.reset
		input  wire        usb_INT1,                   //                  usb.INT1
		inout  wire [15:0] usb_DATA,                   //                     .DATA
		output wire        usb_RST_N,                  //                     .RST_N
		output wire [1:0]  usb_ADDR,                   //                     .ADDR
		output wire        usb_CS_N,                   //                     .CS_N
		output wire        usb_RD_N,                   //                     .RD_N
		output wire        usb_WR_N,                   //                     .WR_N
		input  wire        usb_INT0,                   //                     .INT0
		output wire        vga_CLK,                    //                  vga.CLK
		output wire        vga_HS,                     //                     .HS
		output wire        vga_VS,                     //                     .VS
		output wire        vga_BLANK,                  //                     .BLANK
		output wire        vga_SYNC,                   //                     .SYNC
		output wire [7:0]  vga_R,                      //                     .R
		output wire [7:0]  vga_G,                      //                     .G
		output wire [7:0]  vga_B,                      //                     .B
		input  wire        video_in_TD_CLK27,          //             video_in.TD_CLK27
		input  wire [7:0]  video_in_TD_DATA,           //                     .TD_DATA
		input  wire        video_in_TD_HS,             //                     .TD_HS
		input  wire        video_in_TD_VS,             //                     .TD_VS
		input  wire        video_in_clk27_reset,       //                     .clk27_reset
		output wire        video_in_TD_RESET,          //                     .TD_RESET
		output wire        video_in_overflow_flag,     //                     .overflow_flag
		input  wire        video_pll_ref_clk_clk,      //    video_pll_ref_clk.clk
		input  wire        video_pll_ref_reset_reset   //  video_pll_ref_reset.reset
	);

	wire         system_pll_sys_clk_clk;                                                                // System_PLL:sys_clk_clk -> [AV_Config:clk, Audio_Subsystem:sys_clk_clk, Char_LCD_16x2:clk, Expansion_JP5:clk, Flash:i_clock, Green_LEDs:clk, HEX3_HEX0:clk, HEX7_HEX4:clk, Interval_Timer:clk, Interval_Timer_2:clk, Interval_Timer_2nd_Core:clk, Interval_Timer_2nd_Core_2:clk, IrDA:clk, JTAG_UART:clk, JTAG_UART_2nd_Core:clk, JTAG_to_FPGA_Bridge:clk_clk, Nios2:clk, Nios2_2nd_Core:clk, PS2_Port:clk, PS2_Port_Dual:clk, Pushbuttons:clk, Red_LEDs:clk, SDRAM:clk, SD_Card:i_clock, SRAM:clk, Serial_Port:clk, Slider_Switches:clk, SysID:clock, USB:clk, VGA_Subsystem:sys_clk_clk, Video_In_Subsystem:sys_clk_clk, irq_mapper:clk, irq_mapper_001:clk, mm_interconnect_0:System_PLL_sys_clk_clk, rst_controller:clk, rst_controller_001:clk, rst_controller_002:clk]
	wire         video_pll_vga_clk_clk;                                                                 // Video_PLL:vga_clk_clk -> VGA_Subsystem:vga_clk_clk
	wire         system_pll_reset_source_reset;                                                         // System_PLL:reset_source_reset -> [Audio_Subsystem:sys_reset_reset_n, JTAG_to_FPGA_Bridge:clk_reset_reset, VGA_Subsystem:sys_reset_reset_n, Video_In_Subsystem:sys_reset_reset_n, rst_controller:reset_in0, rst_controller_001:reset_in1, rst_controller_002:reset_in1]
	wire         video_pll_reset_source_reset;                                                          // Video_PLL:reset_source_reset -> VGA_Subsystem:vga_reset_reset_n
	wire  [31:0] nios2_custom_instruction_master_multi_dataa;                                           // Nios2:A_ci_multi_dataa -> Nios2_custom_instruction_master_translator:ci_slave_multi_dataa
	wire         nios2_custom_instruction_master_multi_writerc;                                         // Nios2:A_ci_multi_writerc -> Nios2_custom_instruction_master_translator:ci_slave_multi_writerc
	wire  [31:0] nios2_custom_instruction_master_multi_result;                                          // Nios2_custom_instruction_master_translator:ci_slave_multi_result -> Nios2:A_ci_multi_result
	wire         nios2_custom_instruction_master_clk;                                                   // Nios2:A_ci_multi_clock -> Nios2_custom_instruction_master_translator:ci_slave_multi_clk
	wire  [31:0] nios2_custom_instruction_master_multi_datab;                                           // Nios2:A_ci_multi_datab -> Nios2_custom_instruction_master_translator:ci_slave_multi_datab
	wire         nios2_custom_instruction_master_start;                                                 // Nios2:A_ci_multi_start -> Nios2_custom_instruction_master_translator:ci_slave_multi_start
	wire   [4:0] nios2_custom_instruction_master_multi_b;                                               // Nios2:A_ci_multi_b -> Nios2_custom_instruction_master_translator:ci_slave_multi_b
	wire   [4:0] nios2_custom_instruction_master_multi_c;                                               // Nios2:A_ci_multi_c -> Nios2_custom_instruction_master_translator:ci_slave_multi_c
	wire         nios2_custom_instruction_master_reset_req;                                             // Nios2:A_ci_multi_reset_req -> Nios2_custom_instruction_master_translator:ci_slave_multi_reset_req
	wire         nios2_custom_instruction_master_done;                                                  // Nios2_custom_instruction_master_translator:ci_slave_multi_done -> Nios2:A_ci_multi_done
	wire   [4:0] nios2_custom_instruction_master_multi_a;                                               // Nios2:A_ci_multi_a -> Nios2_custom_instruction_master_translator:ci_slave_multi_a
	wire         nios2_custom_instruction_master_clk_en;                                                // Nios2:A_ci_multi_clk_en -> Nios2_custom_instruction_master_translator:ci_slave_multi_clken
	wire         nios2_custom_instruction_master_reset;                                                 // Nios2:A_ci_multi_reset -> Nios2_custom_instruction_master_translator:ci_slave_multi_reset
	wire         nios2_custom_instruction_master_multi_readrb;                                          // Nios2:A_ci_multi_readrb -> Nios2_custom_instruction_master_translator:ci_slave_multi_readrb
	wire         nios2_custom_instruction_master_multi_readra;                                          // Nios2:A_ci_multi_readra -> Nios2_custom_instruction_master_translator:ci_slave_multi_readra
	wire   [7:0] nios2_custom_instruction_master_multi_n;                                               // Nios2:A_ci_multi_n -> Nios2_custom_instruction_master_translator:ci_slave_multi_n
	wire         nios2_custom_instruction_master_translator_multi_ci_master_readra;                     // Nios2_custom_instruction_master_translator:multi_ci_master_readra -> Nios2_custom_instruction_master_multi_xconnect:ci_slave_readra
	wire   [4:0] nios2_custom_instruction_master_translator_multi_ci_master_a;                          // Nios2_custom_instruction_master_translator:multi_ci_master_a -> Nios2_custom_instruction_master_multi_xconnect:ci_slave_a
	wire   [4:0] nios2_custom_instruction_master_translator_multi_ci_master_b;                          // Nios2_custom_instruction_master_translator:multi_ci_master_b -> Nios2_custom_instruction_master_multi_xconnect:ci_slave_b
	wire         nios2_custom_instruction_master_translator_multi_ci_master_clk;                        // Nios2_custom_instruction_master_translator:multi_ci_master_clk -> Nios2_custom_instruction_master_multi_xconnect:ci_slave_clk
	wire         nios2_custom_instruction_master_translator_multi_ci_master_readrb;                     // Nios2_custom_instruction_master_translator:multi_ci_master_readrb -> Nios2_custom_instruction_master_multi_xconnect:ci_slave_readrb
	wire   [4:0] nios2_custom_instruction_master_translator_multi_ci_master_c;                          // Nios2_custom_instruction_master_translator:multi_ci_master_c -> Nios2_custom_instruction_master_multi_xconnect:ci_slave_c
	wire         nios2_custom_instruction_master_translator_multi_ci_master_start;                      // Nios2_custom_instruction_master_translator:multi_ci_master_start -> Nios2_custom_instruction_master_multi_xconnect:ci_slave_start
	wire         nios2_custom_instruction_master_translator_multi_ci_master_reset_req;                  // Nios2_custom_instruction_master_translator:multi_ci_master_reset_req -> Nios2_custom_instruction_master_multi_xconnect:ci_slave_reset_req
	wire         nios2_custom_instruction_master_translator_multi_ci_master_done;                       // Nios2_custom_instruction_master_multi_xconnect:ci_slave_done -> Nios2_custom_instruction_master_translator:multi_ci_master_done
	wire   [7:0] nios2_custom_instruction_master_translator_multi_ci_master_n;                          // Nios2_custom_instruction_master_translator:multi_ci_master_n -> Nios2_custom_instruction_master_multi_xconnect:ci_slave_n
	wire  [31:0] nios2_custom_instruction_master_translator_multi_ci_master_result;                     // Nios2_custom_instruction_master_multi_xconnect:ci_slave_result -> Nios2_custom_instruction_master_translator:multi_ci_master_result
	wire         nios2_custom_instruction_master_translator_multi_ci_master_clk_en;                     // Nios2_custom_instruction_master_translator:multi_ci_master_clken -> Nios2_custom_instruction_master_multi_xconnect:ci_slave_clken
	wire  [31:0] nios2_custom_instruction_master_translator_multi_ci_master_datab;                      // Nios2_custom_instruction_master_translator:multi_ci_master_datab -> Nios2_custom_instruction_master_multi_xconnect:ci_slave_datab
	wire  [31:0] nios2_custom_instruction_master_translator_multi_ci_master_dataa;                      // Nios2_custom_instruction_master_translator:multi_ci_master_dataa -> Nios2_custom_instruction_master_multi_xconnect:ci_slave_dataa
	wire         nios2_custom_instruction_master_translator_multi_ci_master_reset;                      // Nios2_custom_instruction_master_translator:multi_ci_master_reset -> Nios2_custom_instruction_master_multi_xconnect:ci_slave_reset
	wire         nios2_custom_instruction_master_translator_multi_ci_master_writerc;                    // Nios2_custom_instruction_master_translator:multi_ci_master_writerc -> Nios2_custom_instruction_master_multi_xconnect:ci_slave_writerc
	wire         nios2_custom_instruction_master_multi_xconnect_ci_master0_readra;                      // Nios2_custom_instruction_master_multi_xconnect:ci_master0_readra -> Nios2_custom_instruction_master_multi_slave_translator0:ci_slave_readra
	wire   [4:0] nios2_custom_instruction_master_multi_xconnect_ci_master0_a;                           // Nios2_custom_instruction_master_multi_xconnect:ci_master0_a -> Nios2_custom_instruction_master_multi_slave_translator0:ci_slave_a
	wire   [4:0] nios2_custom_instruction_master_multi_xconnect_ci_master0_b;                           // Nios2_custom_instruction_master_multi_xconnect:ci_master0_b -> Nios2_custom_instruction_master_multi_slave_translator0:ci_slave_b
	wire         nios2_custom_instruction_master_multi_xconnect_ci_master0_readrb;                      // Nios2_custom_instruction_master_multi_xconnect:ci_master0_readrb -> Nios2_custom_instruction_master_multi_slave_translator0:ci_slave_readrb
	wire   [4:0] nios2_custom_instruction_master_multi_xconnect_ci_master0_c;                           // Nios2_custom_instruction_master_multi_xconnect:ci_master0_c -> Nios2_custom_instruction_master_multi_slave_translator0:ci_slave_c
	wire         nios2_custom_instruction_master_multi_xconnect_ci_master0_clk;                         // Nios2_custom_instruction_master_multi_xconnect:ci_master0_clk -> Nios2_custom_instruction_master_multi_slave_translator0:ci_slave_clk
	wire  [31:0] nios2_custom_instruction_master_multi_xconnect_ci_master0_ipending;                    // Nios2_custom_instruction_master_multi_xconnect:ci_master0_ipending -> Nios2_custom_instruction_master_multi_slave_translator0:ci_slave_ipending
	wire         nios2_custom_instruction_master_multi_xconnect_ci_master0_start;                       // Nios2_custom_instruction_master_multi_xconnect:ci_master0_start -> Nios2_custom_instruction_master_multi_slave_translator0:ci_slave_start
	wire         nios2_custom_instruction_master_multi_xconnect_ci_master0_reset_req;                   // Nios2_custom_instruction_master_multi_xconnect:ci_master0_reset_req -> Nios2_custom_instruction_master_multi_slave_translator0:ci_slave_reset_req
	wire         nios2_custom_instruction_master_multi_xconnect_ci_master0_done;                        // Nios2_custom_instruction_master_multi_slave_translator0:ci_slave_done -> Nios2_custom_instruction_master_multi_xconnect:ci_master0_done
	wire   [7:0] nios2_custom_instruction_master_multi_xconnect_ci_master0_n;                           // Nios2_custom_instruction_master_multi_xconnect:ci_master0_n -> Nios2_custom_instruction_master_multi_slave_translator0:ci_slave_n
	wire  [31:0] nios2_custom_instruction_master_multi_xconnect_ci_master0_result;                      // Nios2_custom_instruction_master_multi_slave_translator0:ci_slave_result -> Nios2_custom_instruction_master_multi_xconnect:ci_master0_result
	wire         nios2_custom_instruction_master_multi_xconnect_ci_master0_estatus;                     // Nios2_custom_instruction_master_multi_xconnect:ci_master0_estatus -> Nios2_custom_instruction_master_multi_slave_translator0:ci_slave_estatus
	wire         nios2_custom_instruction_master_multi_xconnect_ci_master0_clk_en;                      // Nios2_custom_instruction_master_multi_xconnect:ci_master0_clken -> Nios2_custom_instruction_master_multi_slave_translator0:ci_slave_clken
	wire  [31:0] nios2_custom_instruction_master_multi_xconnect_ci_master0_datab;                       // Nios2_custom_instruction_master_multi_xconnect:ci_master0_datab -> Nios2_custom_instruction_master_multi_slave_translator0:ci_slave_datab
	wire  [31:0] nios2_custom_instruction_master_multi_xconnect_ci_master0_dataa;                       // Nios2_custom_instruction_master_multi_xconnect:ci_master0_dataa -> Nios2_custom_instruction_master_multi_slave_translator0:ci_slave_dataa
	wire         nios2_custom_instruction_master_multi_xconnect_ci_master0_reset;                       // Nios2_custom_instruction_master_multi_xconnect:ci_master0_reset -> Nios2_custom_instruction_master_multi_slave_translator0:ci_slave_reset
	wire         nios2_custom_instruction_master_multi_xconnect_ci_master0_writerc;                     // Nios2_custom_instruction_master_multi_xconnect:ci_master0_writerc -> Nios2_custom_instruction_master_multi_slave_translator0:ci_slave_writerc
	wire  [31:0] nios2_custom_instruction_master_multi_slave_translator0_ci_master_result;              // Nios2_Floating_Point:result -> Nios2_custom_instruction_master_multi_slave_translator0:ci_master_result
	wire         nios2_custom_instruction_master_multi_slave_translator0_ci_master_clk;                 // Nios2_custom_instruction_master_multi_slave_translator0:ci_master_clk -> Nios2_Floating_Point:clk
	wire         nios2_custom_instruction_master_multi_slave_translator0_ci_master_clk_en;              // Nios2_custom_instruction_master_multi_slave_translator0:ci_master_clken -> Nios2_Floating_Point:clk_en
	wire  [31:0] nios2_custom_instruction_master_multi_slave_translator0_ci_master_datab;               // Nios2_custom_instruction_master_multi_slave_translator0:ci_master_datab -> Nios2_Floating_Point:datab
	wire  [31:0] nios2_custom_instruction_master_multi_slave_translator0_ci_master_dataa;               // Nios2_custom_instruction_master_multi_slave_translator0:ci_master_dataa -> Nios2_Floating_Point:dataa
	wire         nios2_custom_instruction_master_multi_slave_translator0_ci_master_start;               // Nios2_custom_instruction_master_multi_slave_translator0:ci_master_start -> Nios2_Floating_Point:start
	wire         nios2_custom_instruction_master_multi_slave_translator0_ci_master_reset;               // Nios2_custom_instruction_master_multi_slave_translator0:ci_master_reset -> Nios2_Floating_Point:reset
	wire         nios2_custom_instruction_master_multi_slave_translator0_ci_master_done;                // Nios2_Floating_Point:done -> Nios2_custom_instruction_master_multi_slave_translator0:ci_master_done
	wire   [1:0] nios2_custom_instruction_master_multi_slave_translator0_ci_master_n;                   // Nios2_custom_instruction_master_multi_slave_translator0:ci_master_n -> Nios2_Floating_Point:n
	wire         nios2_custom_instruction_master_multi_xconnect_ci_master1_readra;                      // Nios2_custom_instruction_master_multi_xconnect:ci_master1_readra -> Nios2_custom_instruction_master_multi_slave_translator1:ci_slave_readra
	wire   [4:0] nios2_custom_instruction_master_multi_xconnect_ci_master1_a;                           // Nios2_custom_instruction_master_multi_xconnect:ci_master1_a -> Nios2_custom_instruction_master_multi_slave_translator1:ci_slave_a
	wire   [4:0] nios2_custom_instruction_master_multi_xconnect_ci_master1_b;                           // Nios2_custom_instruction_master_multi_xconnect:ci_master1_b -> Nios2_custom_instruction_master_multi_slave_translator1:ci_slave_b
	wire         nios2_custom_instruction_master_multi_xconnect_ci_master1_readrb;                      // Nios2_custom_instruction_master_multi_xconnect:ci_master1_readrb -> Nios2_custom_instruction_master_multi_slave_translator1:ci_slave_readrb
	wire   [4:0] nios2_custom_instruction_master_multi_xconnect_ci_master1_c;                           // Nios2_custom_instruction_master_multi_xconnect:ci_master1_c -> Nios2_custom_instruction_master_multi_slave_translator1:ci_slave_c
	wire         nios2_custom_instruction_master_multi_xconnect_ci_master1_clk;                         // Nios2_custom_instruction_master_multi_xconnect:ci_master1_clk -> Nios2_custom_instruction_master_multi_slave_translator1:ci_slave_clk
	wire  [31:0] nios2_custom_instruction_master_multi_xconnect_ci_master1_ipending;                    // Nios2_custom_instruction_master_multi_xconnect:ci_master1_ipending -> Nios2_custom_instruction_master_multi_slave_translator1:ci_slave_ipending
	wire         nios2_custom_instruction_master_multi_xconnect_ci_master1_start;                       // Nios2_custom_instruction_master_multi_xconnect:ci_master1_start -> Nios2_custom_instruction_master_multi_slave_translator1:ci_slave_start
	wire         nios2_custom_instruction_master_multi_xconnect_ci_master1_reset_req;                   // Nios2_custom_instruction_master_multi_xconnect:ci_master1_reset_req -> Nios2_custom_instruction_master_multi_slave_translator1:ci_slave_reset_req
	wire         nios2_custom_instruction_master_multi_xconnect_ci_master1_done;                        // Nios2_custom_instruction_master_multi_slave_translator1:ci_slave_done -> Nios2_custom_instruction_master_multi_xconnect:ci_master1_done
	wire   [7:0] nios2_custom_instruction_master_multi_xconnect_ci_master1_n;                           // Nios2_custom_instruction_master_multi_xconnect:ci_master1_n -> Nios2_custom_instruction_master_multi_slave_translator1:ci_slave_n
	wire  [31:0] nios2_custom_instruction_master_multi_xconnect_ci_master1_result;                      // Nios2_custom_instruction_master_multi_slave_translator1:ci_slave_result -> Nios2_custom_instruction_master_multi_xconnect:ci_master1_result
	wire         nios2_custom_instruction_master_multi_xconnect_ci_master1_estatus;                     // Nios2_custom_instruction_master_multi_xconnect:ci_master1_estatus -> Nios2_custom_instruction_master_multi_slave_translator1:ci_slave_estatus
	wire         nios2_custom_instruction_master_multi_xconnect_ci_master1_clk_en;                      // Nios2_custom_instruction_master_multi_xconnect:ci_master1_clken -> Nios2_custom_instruction_master_multi_slave_translator1:ci_slave_clken
	wire  [31:0] nios2_custom_instruction_master_multi_xconnect_ci_master1_datab;                       // Nios2_custom_instruction_master_multi_xconnect:ci_master1_datab -> Nios2_custom_instruction_master_multi_slave_translator1:ci_slave_datab
	wire  [31:0] nios2_custom_instruction_master_multi_xconnect_ci_master1_dataa;                       // Nios2_custom_instruction_master_multi_xconnect:ci_master1_dataa -> Nios2_custom_instruction_master_multi_slave_translator1:ci_slave_dataa
	wire         nios2_custom_instruction_master_multi_xconnect_ci_master1_reset;                       // Nios2_custom_instruction_master_multi_xconnect:ci_master1_reset -> Nios2_custom_instruction_master_multi_slave_translator1:ci_slave_reset
	wire         nios2_custom_instruction_master_multi_xconnect_ci_master1_writerc;                     // Nios2_custom_instruction_master_multi_xconnect:ci_master1_writerc -> Nios2_custom_instruction_master_multi_slave_translator1:ci_slave_writerc
	wire  [31:0] nios2_custom_instruction_master_multi_slave_translator1_ci_master_result;              // hw_convolution_inst_0:result -> Nios2_custom_instruction_master_multi_slave_translator1:ci_master_result
	wire         nios2_custom_instruction_master_multi_slave_translator1_ci_master_clk;                 // Nios2_custom_instruction_master_multi_slave_translator1:ci_master_clk -> hw_convolution_inst_0:clk
	wire         nios2_custom_instruction_master_multi_slave_translator1_ci_master_clk_en;              // Nios2_custom_instruction_master_multi_slave_translator1:ci_master_clken -> hw_convolution_inst_0:clk_en
	wire  [31:0] nios2_custom_instruction_master_multi_slave_translator1_ci_master_datab;               // Nios2_custom_instruction_master_multi_slave_translator1:ci_master_datab -> hw_convolution_inst_0:datab
	wire  [31:0] nios2_custom_instruction_master_multi_slave_translator1_ci_master_dataa;               // Nios2_custom_instruction_master_multi_slave_translator1:ci_master_dataa -> hw_convolution_inst_0:dataa
	wire         nios2_custom_instruction_master_multi_slave_translator1_ci_master_start;               // Nios2_custom_instruction_master_multi_slave_translator1:ci_master_start -> hw_convolution_inst_0:start
	wire         nios2_custom_instruction_master_multi_slave_translator1_ci_master_reset;               // Nios2_custom_instruction_master_multi_slave_translator1:ci_master_reset -> hw_convolution_inst_0:reset
	wire         nios2_custom_instruction_master_multi_slave_translator1_ci_master_done;                // hw_convolution_inst_0:done -> Nios2_custom_instruction_master_multi_slave_translator1:ci_master_done
	wire  [31:0] nios2_2nd_core_custom_instruction_master_multi_dataa;                                  // Nios2_2nd_Core:A_ci_multi_dataa -> Nios2_2nd_Core_custom_instruction_master_translator:ci_slave_multi_dataa
	wire         nios2_2nd_core_custom_instruction_master_multi_writerc;                                // Nios2_2nd_Core:A_ci_multi_writerc -> Nios2_2nd_Core_custom_instruction_master_translator:ci_slave_multi_writerc
	wire  [31:0] nios2_2nd_core_custom_instruction_master_multi_result;                                 // Nios2_2nd_Core_custom_instruction_master_translator:ci_slave_multi_result -> Nios2_2nd_Core:A_ci_multi_result
	wire         nios2_2nd_core_custom_instruction_master_clk;                                          // Nios2_2nd_Core:A_ci_multi_clock -> Nios2_2nd_Core_custom_instruction_master_translator:ci_slave_multi_clk
	wire  [31:0] nios2_2nd_core_custom_instruction_master_multi_datab;                                  // Nios2_2nd_Core:A_ci_multi_datab -> Nios2_2nd_Core_custom_instruction_master_translator:ci_slave_multi_datab
	wire         nios2_2nd_core_custom_instruction_master_start;                                        // Nios2_2nd_Core:A_ci_multi_start -> Nios2_2nd_Core_custom_instruction_master_translator:ci_slave_multi_start
	wire   [4:0] nios2_2nd_core_custom_instruction_master_multi_b;                                      // Nios2_2nd_Core:A_ci_multi_b -> Nios2_2nd_Core_custom_instruction_master_translator:ci_slave_multi_b
	wire   [4:0] nios2_2nd_core_custom_instruction_master_multi_c;                                      // Nios2_2nd_Core:A_ci_multi_c -> Nios2_2nd_Core_custom_instruction_master_translator:ci_slave_multi_c
	wire         nios2_2nd_core_custom_instruction_master_reset_req;                                    // Nios2_2nd_Core:A_ci_multi_reset_req -> Nios2_2nd_Core_custom_instruction_master_translator:ci_slave_multi_reset_req
	wire         nios2_2nd_core_custom_instruction_master_done;                                         // Nios2_2nd_Core_custom_instruction_master_translator:ci_slave_multi_done -> Nios2_2nd_Core:A_ci_multi_done
	wire   [4:0] nios2_2nd_core_custom_instruction_master_multi_a;                                      // Nios2_2nd_Core:A_ci_multi_a -> Nios2_2nd_Core_custom_instruction_master_translator:ci_slave_multi_a
	wire         nios2_2nd_core_custom_instruction_master_clk_en;                                       // Nios2_2nd_Core:A_ci_multi_clk_en -> Nios2_2nd_Core_custom_instruction_master_translator:ci_slave_multi_clken
	wire         nios2_2nd_core_custom_instruction_master_reset;                                        // Nios2_2nd_Core:A_ci_multi_reset -> Nios2_2nd_Core_custom_instruction_master_translator:ci_slave_multi_reset
	wire         nios2_2nd_core_custom_instruction_master_multi_readrb;                                 // Nios2_2nd_Core:A_ci_multi_readrb -> Nios2_2nd_Core_custom_instruction_master_translator:ci_slave_multi_readrb
	wire         nios2_2nd_core_custom_instruction_master_multi_readra;                                 // Nios2_2nd_Core:A_ci_multi_readra -> Nios2_2nd_Core_custom_instruction_master_translator:ci_slave_multi_readra
	wire   [7:0] nios2_2nd_core_custom_instruction_master_multi_n;                                      // Nios2_2nd_Core:A_ci_multi_n -> Nios2_2nd_Core_custom_instruction_master_translator:ci_slave_multi_n
	wire         nios2_2nd_core_custom_instruction_master_translator_multi_ci_master_readra;            // Nios2_2nd_Core_custom_instruction_master_translator:multi_ci_master_readra -> Nios2_2nd_Core_custom_instruction_master_multi_xconnect:ci_slave_readra
	wire   [4:0] nios2_2nd_core_custom_instruction_master_translator_multi_ci_master_a;                 // Nios2_2nd_Core_custom_instruction_master_translator:multi_ci_master_a -> Nios2_2nd_Core_custom_instruction_master_multi_xconnect:ci_slave_a
	wire   [4:0] nios2_2nd_core_custom_instruction_master_translator_multi_ci_master_b;                 // Nios2_2nd_Core_custom_instruction_master_translator:multi_ci_master_b -> Nios2_2nd_Core_custom_instruction_master_multi_xconnect:ci_slave_b
	wire         nios2_2nd_core_custom_instruction_master_translator_multi_ci_master_clk;               // Nios2_2nd_Core_custom_instruction_master_translator:multi_ci_master_clk -> Nios2_2nd_Core_custom_instruction_master_multi_xconnect:ci_slave_clk
	wire         nios2_2nd_core_custom_instruction_master_translator_multi_ci_master_readrb;            // Nios2_2nd_Core_custom_instruction_master_translator:multi_ci_master_readrb -> Nios2_2nd_Core_custom_instruction_master_multi_xconnect:ci_slave_readrb
	wire   [4:0] nios2_2nd_core_custom_instruction_master_translator_multi_ci_master_c;                 // Nios2_2nd_Core_custom_instruction_master_translator:multi_ci_master_c -> Nios2_2nd_Core_custom_instruction_master_multi_xconnect:ci_slave_c
	wire         nios2_2nd_core_custom_instruction_master_translator_multi_ci_master_start;             // Nios2_2nd_Core_custom_instruction_master_translator:multi_ci_master_start -> Nios2_2nd_Core_custom_instruction_master_multi_xconnect:ci_slave_start
	wire         nios2_2nd_core_custom_instruction_master_translator_multi_ci_master_reset_req;         // Nios2_2nd_Core_custom_instruction_master_translator:multi_ci_master_reset_req -> Nios2_2nd_Core_custom_instruction_master_multi_xconnect:ci_slave_reset_req
	wire         nios2_2nd_core_custom_instruction_master_translator_multi_ci_master_done;              // Nios2_2nd_Core_custom_instruction_master_multi_xconnect:ci_slave_done -> Nios2_2nd_Core_custom_instruction_master_translator:multi_ci_master_done
	wire   [7:0] nios2_2nd_core_custom_instruction_master_translator_multi_ci_master_n;                 // Nios2_2nd_Core_custom_instruction_master_translator:multi_ci_master_n -> Nios2_2nd_Core_custom_instruction_master_multi_xconnect:ci_slave_n
	wire  [31:0] nios2_2nd_core_custom_instruction_master_translator_multi_ci_master_result;            // Nios2_2nd_Core_custom_instruction_master_multi_xconnect:ci_slave_result -> Nios2_2nd_Core_custom_instruction_master_translator:multi_ci_master_result
	wire         nios2_2nd_core_custom_instruction_master_translator_multi_ci_master_clk_en;            // Nios2_2nd_Core_custom_instruction_master_translator:multi_ci_master_clken -> Nios2_2nd_Core_custom_instruction_master_multi_xconnect:ci_slave_clken
	wire  [31:0] nios2_2nd_core_custom_instruction_master_translator_multi_ci_master_datab;             // Nios2_2nd_Core_custom_instruction_master_translator:multi_ci_master_datab -> Nios2_2nd_Core_custom_instruction_master_multi_xconnect:ci_slave_datab
	wire  [31:0] nios2_2nd_core_custom_instruction_master_translator_multi_ci_master_dataa;             // Nios2_2nd_Core_custom_instruction_master_translator:multi_ci_master_dataa -> Nios2_2nd_Core_custom_instruction_master_multi_xconnect:ci_slave_dataa
	wire         nios2_2nd_core_custom_instruction_master_translator_multi_ci_master_reset;             // Nios2_2nd_Core_custom_instruction_master_translator:multi_ci_master_reset -> Nios2_2nd_Core_custom_instruction_master_multi_xconnect:ci_slave_reset
	wire         nios2_2nd_core_custom_instruction_master_translator_multi_ci_master_writerc;           // Nios2_2nd_Core_custom_instruction_master_translator:multi_ci_master_writerc -> Nios2_2nd_Core_custom_instruction_master_multi_xconnect:ci_slave_writerc
	wire         nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_readra;             // Nios2_2nd_Core_custom_instruction_master_multi_xconnect:ci_master0_readra -> Nios2_2nd_Core_custom_instruction_master_multi_slave_translator0:ci_slave_readra
	wire   [4:0] nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_a;                  // Nios2_2nd_Core_custom_instruction_master_multi_xconnect:ci_master0_a -> Nios2_2nd_Core_custom_instruction_master_multi_slave_translator0:ci_slave_a
	wire   [4:0] nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_b;                  // Nios2_2nd_Core_custom_instruction_master_multi_xconnect:ci_master0_b -> Nios2_2nd_Core_custom_instruction_master_multi_slave_translator0:ci_slave_b
	wire         nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_readrb;             // Nios2_2nd_Core_custom_instruction_master_multi_xconnect:ci_master0_readrb -> Nios2_2nd_Core_custom_instruction_master_multi_slave_translator0:ci_slave_readrb
	wire   [4:0] nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_c;                  // Nios2_2nd_Core_custom_instruction_master_multi_xconnect:ci_master0_c -> Nios2_2nd_Core_custom_instruction_master_multi_slave_translator0:ci_slave_c
	wire         nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_clk;                // Nios2_2nd_Core_custom_instruction_master_multi_xconnect:ci_master0_clk -> Nios2_2nd_Core_custom_instruction_master_multi_slave_translator0:ci_slave_clk
	wire  [31:0] nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_ipending;           // Nios2_2nd_Core_custom_instruction_master_multi_xconnect:ci_master0_ipending -> Nios2_2nd_Core_custom_instruction_master_multi_slave_translator0:ci_slave_ipending
	wire         nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_start;              // Nios2_2nd_Core_custom_instruction_master_multi_xconnect:ci_master0_start -> Nios2_2nd_Core_custom_instruction_master_multi_slave_translator0:ci_slave_start
	wire         nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_reset_req;          // Nios2_2nd_Core_custom_instruction_master_multi_xconnect:ci_master0_reset_req -> Nios2_2nd_Core_custom_instruction_master_multi_slave_translator0:ci_slave_reset_req
	wire         nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_done;               // Nios2_2nd_Core_custom_instruction_master_multi_slave_translator0:ci_slave_done -> Nios2_2nd_Core_custom_instruction_master_multi_xconnect:ci_master0_done
	wire   [7:0] nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_n;                  // Nios2_2nd_Core_custom_instruction_master_multi_xconnect:ci_master0_n -> Nios2_2nd_Core_custom_instruction_master_multi_slave_translator0:ci_slave_n
	wire  [31:0] nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_result;             // Nios2_2nd_Core_custom_instruction_master_multi_slave_translator0:ci_slave_result -> Nios2_2nd_Core_custom_instruction_master_multi_xconnect:ci_master0_result
	wire         nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_estatus;            // Nios2_2nd_Core_custom_instruction_master_multi_xconnect:ci_master0_estatus -> Nios2_2nd_Core_custom_instruction_master_multi_slave_translator0:ci_slave_estatus
	wire         nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_clk_en;             // Nios2_2nd_Core_custom_instruction_master_multi_xconnect:ci_master0_clken -> Nios2_2nd_Core_custom_instruction_master_multi_slave_translator0:ci_slave_clken
	wire  [31:0] nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_datab;              // Nios2_2nd_Core_custom_instruction_master_multi_xconnect:ci_master0_datab -> Nios2_2nd_Core_custom_instruction_master_multi_slave_translator0:ci_slave_datab
	wire  [31:0] nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_dataa;              // Nios2_2nd_Core_custom_instruction_master_multi_xconnect:ci_master0_dataa -> Nios2_2nd_Core_custom_instruction_master_multi_slave_translator0:ci_slave_dataa
	wire         nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_reset;              // Nios2_2nd_Core_custom_instruction_master_multi_xconnect:ci_master0_reset -> Nios2_2nd_Core_custom_instruction_master_multi_slave_translator0:ci_slave_reset
	wire         nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_writerc;            // Nios2_2nd_Core_custom_instruction_master_multi_xconnect:ci_master0_writerc -> Nios2_2nd_Core_custom_instruction_master_multi_slave_translator0:ci_slave_writerc
	wire  [31:0] nios2_2nd_core_custom_instruction_master_multi_slave_translator0_ci_master_result;     // Nios2_2nd_Core_Floating_Point:result -> Nios2_2nd_Core_custom_instruction_master_multi_slave_translator0:ci_master_result
	wire         nios2_2nd_core_custom_instruction_master_multi_slave_translator0_ci_master_clk;        // Nios2_2nd_Core_custom_instruction_master_multi_slave_translator0:ci_master_clk -> Nios2_2nd_Core_Floating_Point:clk
	wire         nios2_2nd_core_custom_instruction_master_multi_slave_translator0_ci_master_clk_en;     // Nios2_2nd_Core_custom_instruction_master_multi_slave_translator0:ci_master_clken -> Nios2_2nd_Core_Floating_Point:clk_en
	wire  [31:0] nios2_2nd_core_custom_instruction_master_multi_slave_translator0_ci_master_datab;      // Nios2_2nd_Core_custom_instruction_master_multi_slave_translator0:ci_master_datab -> Nios2_2nd_Core_Floating_Point:datab
	wire  [31:0] nios2_2nd_core_custom_instruction_master_multi_slave_translator0_ci_master_dataa;      // Nios2_2nd_Core_custom_instruction_master_multi_slave_translator0:ci_master_dataa -> Nios2_2nd_Core_Floating_Point:dataa
	wire         nios2_2nd_core_custom_instruction_master_multi_slave_translator0_ci_master_start;      // Nios2_2nd_Core_custom_instruction_master_multi_slave_translator0:ci_master_start -> Nios2_2nd_Core_Floating_Point:start
	wire         nios2_2nd_core_custom_instruction_master_multi_slave_translator0_ci_master_reset;      // Nios2_2nd_Core_custom_instruction_master_multi_slave_translator0:ci_master_reset -> Nios2_2nd_Core_Floating_Point:reset
	wire         nios2_2nd_core_custom_instruction_master_multi_slave_translator0_ci_master_done;       // Nios2_2nd_Core_Floating_Point:done -> Nios2_2nd_Core_custom_instruction_master_multi_slave_translator0:ci_master_done
	wire   [1:0] nios2_2nd_core_custom_instruction_master_multi_slave_translator0_ci_master_n;          // Nios2_2nd_Core_custom_instruction_master_multi_slave_translator0:ci_master_n -> Nios2_2nd_Core_Floating_Point:n
	wire  [31:0] nios2_data_master_readdata;                                                            // mm_interconnect_0:Nios2_data_master_readdata -> Nios2:d_readdata
	wire         nios2_data_master_waitrequest;                                                         // mm_interconnect_0:Nios2_data_master_waitrequest -> Nios2:d_waitrequest
	wire         nios2_data_master_debugaccess;                                                         // Nios2:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:Nios2_data_master_debugaccess
	wire  [31:0] nios2_data_master_address;                                                             // Nios2:d_address -> mm_interconnect_0:Nios2_data_master_address
	wire   [3:0] nios2_data_master_byteenable;                                                          // Nios2:d_byteenable -> mm_interconnect_0:Nios2_data_master_byteenable
	wire         nios2_data_master_read;                                                                // Nios2:d_read -> mm_interconnect_0:Nios2_data_master_read
	wire         nios2_data_master_write;                                                               // Nios2:d_write -> mm_interconnect_0:Nios2_data_master_write
	wire  [31:0] nios2_data_master_writedata;                                                           // Nios2:d_writedata -> mm_interconnect_0:Nios2_data_master_writedata
	wire  [31:0] nios2_2nd_core_data_master_readdata;                                                   // mm_interconnect_0:Nios2_2nd_Core_data_master_readdata -> Nios2_2nd_Core:d_readdata
	wire         nios2_2nd_core_data_master_waitrequest;                                                // mm_interconnect_0:Nios2_2nd_Core_data_master_waitrequest -> Nios2_2nd_Core:d_waitrequest
	wire         nios2_2nd_core_data_master_debugaccess;                                                // Nios2_2nd_Core:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:Nios2_2nd_Core_data_master_debugaccess
	wire  [31:0] nios2_2nd_core_data_master_address;                                                    // Nios2_2nd_Core:d_address -> mm_interconnect_0:Nios2_2nd_Core_data_master_address
	wire   [3:0] nios2_2nd_core_data_master_byteenable;                                                 // Nios2_2nd_Core:d_byteenable -> mm_interconnect_0:Nios2_2nd_Core_data_master_byteenable
	wire         nios2_2nd_core_data_master_read;                                                       // Nios2_2nd_Core:d_read -> mm_interconnect_0:Nios2_2nd_Core_data_master_read
	wire         nios2_2nd_core_data_master_write;                                                      // Nios2_2nd_Core:d_write -> mm_interconnect_0:Nios2_2nd_Core_data_master_write
	wire  [31:0] nios2_2nd_core_data_master_writedata;                                                  // Nios2_2nd_Core:d_writedata -> mm_interconnect_0:Nios2_2nd_Core_data_master_writedata
	wire  [31:0] jtag_to_fpga_bridge_master_readdata;                                                   // mm_interconnect_0:JTAG_to_FPGA_Bridge_master_readdata -> JTAG_to_FPGA_Bridge:master_readdata
	wire         jtag_to_fpga_bridge_master_waitrequest;                                                // mm_interconnect_0:JTAG_to_FPGA_Bridge_master_waitrequest -> JTAG_to_FPGA_Bridge:master_waitrequest
	wire  [31:0] jtag_to_fpga_bridge_master_address;                                                    // JTAG_to_FPGA_Bridge:master_address -> mm_interconnect_0:JTAG_to_FPGA_Bridge_master_address
	wire         jtag_to_fpga_bridge_master_read;                                                       // JTAG_to_FPGA_Bridge:master_read -> mm_interconnect_0:JTAG_to_FPGA_Bridge_master_read
	wire   [3:0] jtag_to_fpga_bridge_master_byteenable;                                                 // JTAG_to_FPGA_Bridge:master_byteenable -> mm_interconnect_0:JTAG_to_FPGA_Bridge_master_byteenable
	wire         jtag_to_fpga_bridge_master_readdatavalid;                                              // mm_interconnect_0:JTAG_to_FPGA_Bridge_master_readdatavalid -> JTAG_to_FPGA_Bridge:master_readdatavalid
	wire         jtag_to_fpga_bridge_master_write;                                                      // JTAG_to_FPGA_Bridge:master_write -> mm_interconnect_0:JTAG_to_FPGA_Bridge_master_write
	wire  [31:0] jtag_to_fpga_bridge_master_writedata;                                                  // JTAG_to_FPGA_Bridge:master_writedata -> mm_interconnect_0:JTAG_to_FPGA_Bridge_master_writedata
	wire  [31:0] nios2_2nd_core_instruction_master_readdata;                                            // mm_interconnect_0:Nios2_2nd_Core_instruction_master_readdata -> Nios2_2nd_Core:i_readdata
	wire         nios2_2nd_core_instruction_master_waitrequest;                                         // mm_interconnect_0:Nios2_2nd_Core_instruction_master_waitrequest -> Nios2_2nd_Core:i_waitrequest
	wire  [27:0] nios2_2nd_core_instruction_master_address;                                             // Nios2_2nd_Core:i_address -> mm_interconnect_0:Nios2_2nd_Core_instruction_master_address
	wire         nios2_2nd_core_instruction_master_read;                                                // Nios2_2nd_Core:i_read -> mm_interconnect_0:Nios2_2nd_Core_instruction_master_read
	wire         nios2_2nd_core_instruction_master_readdatavalid;                                       // mm_interconnect_0:Nios2_2nd_Core_instruction_master_readdatavalid -> Nios2_2nd_Core:i_readdatavalid
	wire  [31:0] nios2_instruction_master_readdata;                                                     // mm_interconnect_0:Nios2_instruction_master_readdata -> Nios2:i_readdata
	wire         nios2_instruction_master_waitrequest;                                                  // mm_interconnect_0:Nios2_instruction_master_waitrequest -> Nios2:i_waitrequest
	wire  [27:0] nios2_instruction_master_address;                                                      // Nios2:i_address -> mm_interconnect_0:Nios2_instruction_master_address
	wire         nios2_instruction_master_read;                                                         // Nios2:i_read -> mm_interconnect_0:Nios2_instruction_master_read
	wire         nios2_instruction_master_readdatavalid;                                                // mm_interconnect_0:Nios2_instruction_master_readdatavalid -> Nios2:i_readdatavalid
	wire         vga_subsystem_pixel_dma_master_waitrequest;                                            // mm_interconnect_0:VGA_Subsystem_pixel_dma_master_waitrequest -> VGA_Subsystem:pixel_dma_master_waitrequest
	wire  [15:0] vga_subsystem_pixel_dma_master_readdata;                                               // mm_interconnect_0:VGA_Subsystem_pixel_dma_master_readdata -> VGA_Subsystem:pixel_dma_master_readdata
	wire  [31:0] vga_subsystem_pixel_dma_master_address;                                                // VGA_Subsystem:pixel_dma_master_address -> mm_interconnect_0:VGA_Subsystem_pixel_dma_master_address
	wire         vga_subsystem_pixel_dma_master_read;                                                   // VGA_Subsystem:pixel_dma_master_read -> mm_interconnect_0:VGA_Subsystem_pixel_dma_master_read
	wire         vga_subsystem_pixel_dma_master_readdatavalid;                                          // mm_interconnect_0:VGA_Subsystem_pixel_dma_master_readdatavalid -> VGA_Subsystem:pixel_dma_master_readdatavalid
	wire         vga_subsystem_pixel_dma_master_lock;                                                   // VGA_Subsystem:pixel_dma_master_lock -> mm_interconnect_0:VGA_Subsystem_pixel_dma_master_lock
	wire         video_in_subsystem_video_in_dma_master_waitrequest;                                    // mm_interconnect_0:Video_In_Subsystem_video_in_dma_master_waitrequest -> Video_In_Subsystem:video_in_dma_master_waitrequest
	wire  [31:0] video_in_subsystem_video_in_dma_master_address;                                        // Video_In_Subsystem:video_in_dma_master_address -> mm_interconnect_0:Video_In_Subsystem_video_in_dma_master_address
	wire         video_in_subsystem_video_in_dma_master_write;                                          // Video_In_Subsystem:video_in_dma_master_write -> mm_interconnect_0:Video_In_Subsystem_video_in_dma_master_write
	wire  [15:0] video_in_subsystem_video_in_dma_master_writedata;                                      // Video_In_Subsystem:video_in_dma_master_writedata -> mm_interconnect_0:Video_In_Subsystem_video_in_dma_master_writedata
	wire         mm_interconnect_0_audio_subsystem_audio_slave_chipselect;                              // mm_interconnect_0:Audio_Subsystem_audio_slave_chipselect -> Audio_Subsystem:audio_slave_chipselect
	wire  [31:0] mm_interconnect_0_audio_subsystem_audio_slave_readdata;                                // Audio_Subsystem:audio_slave_readdata -> mm_interconnect_0:Audio_Subsystem_audio_slave_readdata
	wire   [1:0] mm_interconnect_0_audio_subsystem_audio_slave_address;                                 // mm_interconnect_0:Audio_Subsystem_audio_slave_address -> Audio_Subsystem:audio_slave_address
	wire         mm_interconnect_0_audio_subsystem_audio_slave_read;                                    // mm_interconnect_0:Audio_Subsystem_audio_slave_read -> Audio_Subsystem:audio_slave_read
	wire         mm_interconnect_0_audio_subsystem_audio_slave_write;                                   // mm_interconnect_0:Audio_Subsystem_audio_slave_write -> Audio_Subsystem:audio_slave_write
	wire  [31:0] mm_interconnect_0_audio_subsystem_audio_slave_writedata;                               // mm_interconnect_0:Audio_Subsystem_audio_slave_writedata -> Audio_Subsystem:audio_slave_writedata
	wire  [31:0] mm_interconnect_0_av_config_avalon_av_config_slave_readdata;                           // AV_Config:readdata -> mm_interconnect_0:AV_Config_avalon_av_config_slave_readdata
	wire         mm_interconnect_0_av_config_avalon_av_config_slave_waitrequest;                        // AV_Config:waitrequest -> mm_interconnect_0:AV_Config_avalon_av_config_slave_waitrequest
	wire   [1:0] mm_interconnect_0_av_config_avalon_av_config_slave_address;                            // mm_interconnect_0:AV_Config_avalon_av_config_slave_address -> AV_Config:address
	wire         mm_interconnect_0_av_config_avalon_av_config_slave_read;                               // mm_interconnect_0:AV_Config_avalon_av_config_slave_read -> AV_Config:read
	wire   [3:0] mm_interconnect_0_av_config_avalon_av_config_slave_byteenable;                         // mm_interconnect_0:AV_Config_avalon_av_config_slave_byteenable -> AV_Config:byteenable
	wire         mm_interconnect_0_av_config_avalon_av_config_slave_write;                              // mm_interconnect_0:AV_Config_avalon_av_config_slave_write -> AV_Config:write
	wire  [31:0] mm_interconnect_0_av_config_avalon_av_config_slave_writedata;                          // mm_interconnect_0:AV_Config_avalon_av_config_slave_writedata -> AV_Config:writedata
	wire         mm_interconnect_0_irda_avalon_irda_slave_chipselect;                                   // mm_interconnect_0:IrDA_avalon_irda_slave_chipselect -> IrDA:chipselect
	wire  [31:0] mm_interconnect_0_irda_avalon_irda_slave_readdata;                                     // IrDA:readdata -> mm_interconnect_0:IrDA_avalon_irda_slave_readdata
	wire   [0:0] mm_interconnect_0_irda_avalon_irda_slave_address;                                      // mm_interconnect_0:IrDA_avalon_irda_slave_address -> IrDA:address
	wire         mm_interconnect_0_irda_avalon_irda_slave_read;                                         // mm_interconnect_0:IrDA_avalon_irda_slave_read -> IrDA:read
	wire   [3:0] mm_interconnect_0_irda_avalon_irda_slave_byteenable;                                   // mm_interconnect_0:IrDA_avalon_irda_slave_byteenable -> IrDA:byteenable
	wire         mm_interconnect_0_irda_avalon_irda_slave_write;                                        // mm_interconnect_0:IrDA_avalon_irda_slave_write -> IrDA:write
	wire  [31:0] mm_interconnect_0_irda_avalon_irda_slave_writedata;                                    // mm_interconnect_0:IrDA_avalon_irda_slave_writedata -> IrDA:writedata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;                              // mm_interconnect_0:JTAG_UART_avalon_jtag_slave_chipselect -> JTAG_UART:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;                                // JTAG_UART:av_readdata -> mm_interconnect_0:JTAG_UART_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest;                             // JTAG_UART:av_waitrequest -> mm_interconnect_0:JTAG_UART_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;                                 // mm_interconnect_0:JTAG_UART_avalon_jtag_slave_address -> JTAG_UART:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;                                    // mm_interconnect_0:JTAG_UART_avalon_jtag_slave_read -> JTAG_UART:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;                                   // mm_interconnect_0:JTAG_UART_avalon_jtag_slave_write -> JTAG_UART:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;                               // mm_interconnect_0:JTAG_UART_avalon_jtag_slave_writedata -> JTAG_UART:av_writedata
	wire         mm_interconnect_0_char_lcd_16x2_avalon_lcd_slave_chipselect;                           // mm_interconnect_0:Char_LCD_16x2_avalon_lcd_slave_chipselect -> Char_LCD_16x2:chipselect
	wire   [7:0] mm_interconnect_0_char_lcd_16x2_avalon_lcd_slave_readdata;                             // Char_LCD_16x2:readdata -> mm_interconnect_0:Char_LCD_16x2_avalon_lcd_slave_readdata
	wire         mm_interconnect_0_char_lcd_16x2_avalon_lcd_slave_waitrequest;                          // Char_LCD_16x2:waitrequest -> mm_interconnect_0:Char_LCD_16x2_avalon_lcd_slave_waitrequest
	wire   [0:0] mm_interconnect_0_char_lcd_16x2_avalon_lcd_slave_address;                              // mm_interconnect_0:Char_LCD_16x2_avalon_lcd_slave_address -> Char_LCD_16x2:address
	wire         mm_interconnect_0_char_lcd_16x2_avalon_lcd_slave_read;                                 // mm_interconnect_0:Char_LCD_16x2_avalon_lcd_slave_read -> Char_LCD_16x2:read
	wire         mm_interconnect_0_char_lcd_16x2_avalon_lcd_slave_write;                                // mm_interconnect_0:Char_LCD_16x2_avalon_lcd_slave_write -> Char_LCD_16x2:write
	wire   [7:0] mm_interconnect_0_char_lcd_16x2_avalon_lcd_slave_writedata;                            // mm_interconnect_0:Char_LCD_16x2_avalon_lcd_slave_writedata -> Char_LCD_16x2:writedata
	wire         mm_interconnect_0_ps2_port_avalon_ps2_slave_chipselect;                                // mm_interconnect_0:PS2_Port_avalon_ps2_slave_chipselect -> PS2_Port:chipselect
	wire  [31:0] mm_interconnect_0_ps2_port_avalon_ps2_slave_readdata;                                  // PS2_Port:readdata -> mm_interconnect_0:PS2_Port_avalon_ps2_slave_readdata
	wire         mm_interconnect_0_ps2_port_avalon_ps2_slave_waitrequest;                               // PS2_Port:waitrequest -> mm_interconnect_0:PS2_Port_avalon_ps2_slave_waitrequest
	wire   [0:0] mm_interconnect_0_ps2_port_avalon_ps2_slave_address;                                   // mm_interconnect_0:PS2_Port_avalon_ps2_slave_address -> PS2_Port:address
	wire         mm_interconnect_0_ps2_port_avalon_ps2_slave_read;                                      // mm_interconnect_0:PS2_Port_avalon_ps2_slave_read -> PS2_Port:read
	wire   [3:0] mm_interconnect_0_ps2_port_avalon_ps2_slave_byteenable;                                // mm_interconnect_0:PS2_Port_avalon_ps2_slave_byteenable -> PS2_Port:byteenable
	wire         mm_interconnect_0_ps2_port_avalon_ps2_slave_write;                                     // mm_interconnect_0:PS2_Port_avalon_ps2_slave_write -> PS2_Port:write
	wire  [31:0] mm_interconnect_0_ps2_port_avalon_ps2_slave_writedata;                                 // mm_interconnect_0:PS2_Port_avalon_ps2_slave_writedata -> PS2_Port:writedata
	wire         mm_interconnect_0_ps2_port_dual_avalon_ps2_slave_chipselect;                           // mm_interconnect_0:PS2_Port_Dual_avalon_ps2_slave_chipselect -> PS2_Port_Dual:chipselect
	wire  [31:0] mm_interconnect_0_ps2_port_dual_avalon_ps2_slave_readdata;                             // PS2_Port_Dual:readdata -> mm_interconnect_0:PS2_Port_Dual_avalon_ps2_slave_readdata
	wire         mm_interconnect_0_ps2_port_dual_avalon_ps2_slave_waitrequest;                          // PS2_Port_Dual:waitrequest -> mm_interconnect_0:PS2_Port_Dual_avalon_ps2_slave_waitrequest
	wire   [0:0] mm_interconnect_0_ps2_port_dual_avalon_ps2_slave_address;                              // mm_interconnect_0:PS2_Port_Dual_avalon_ps2_slave_address -> PS2_Port_Dual:address
	wire         mm_interconnect_0_ps2_port_dual_avalon_ps2_slave_read;                                 // mm_interconnect_0:PS2_Port_Dual_avalon_ps2_slave_read -> PS2_Port_Dual:read
	wire   [3:0] mm_interconnect_0_ps2_port_dual_avalon_ps2_slave_byteenable;                           // mm_interconnect_0:PS2_Port_Dual_avalon_ps2_slave_byteenable -> PS2_Port_Dual:byteenable
	wire         mm_interconnect_0_ps2_port_dual_avalon_ps2_slave_write;                                // mm_interconnect_0:PS2_Port_Dual_avalon_ps2_slave_write -> PS2_Port_Dual:write
	wire  [31:0] mm_interconnect_0_ps2_port_dual_avalon_ps2_slave_writedata;                            // mm_interconnect_0:PS2_Port_Dual_avalon_ps2_slave_writedata -> PS2_Port_Dual:writedata
	wire         mm_interconnect_0_serial_port_avalon_rs232_slave_chipselect;                           // mm_interconnect_0:Serial_Port_avalon_rs232_slave_chipselect -> Serial_Port:chipselect
	wire  [31:0] mm_interconnect_0_serial_port_avalon_rs232_slave_readdata;                             // Serial_Port:readdata -> mm_interconnect_0:Serial_Port_avalon_rs232_slave_readdata
	wire   [0:0] mm_interconnect_0_serial_port_avalon_rs232_slave_address;                              // mm_interconnect_0:Serial_Port_avalon_rs232_slave_address -> Serial_Port:address
	wire         mm_interconnect_0_serial_port_avalon_rs232_slave_read;                                 // mm_interconnect_0:Serial_Port_avalon_rs232_slave_read -> Serial_Port:read
	wire   [3:0] mm_interconnect_0_serial_port_avalon_rs232_slave_byteenable;                           // mm_interconnect_0:Serial_Port_avalon_rs232_slave_byteenable -> Serial_Port:byteenable
	wire         mm_interconnect_0_serial_port_avalon_rs232_slave_write;                                // mm_interconnect_0:Serial_Port_avalon_rs232_slave_write -> Serial_Port:write
	wire  [31:0] mm_interconnect_0_serial_port_avalon_rs232_slave_writedata;                            // mm_interconnect_0:Serial_Port_avalon_rs232_slave_writedata -> Serial_Port:writedata
	wire         mm_interconnect_0_sd_card_avalon_sdcard_slave_chipselect;                              // mm_interconnect_0:SD_Card_avalon_sdcard_slave_chipselect -> SD_Card:i_avalon_chip_select
	wire  [31:0] mm_interconnect_0_sd_card_avalon_sdcard_slave_readdata;                                // SD_Card:o_avalon_readdata -> mm_interconnect_0:SD_Card_avalon_sdcard_slave_readdata
	wire         mm_interconnect_0_sd_card_avalon_sdcard_slave_waitrequest;                             // SD_Card:o_avalon_waitrequest -> mm_interconnect_0:SD_Card_avalon_sdcard_slave_waitrequest
	wire   [7:0] mm_interconnect_0_sd_card_avalon_sdcard_slave_address;                                 // mm_interconnect_0:SD_Card_avalon_sdcard_slave_address -> SD_Card:i_avalon_address
	wire         mm_interconnect_0_sd_card_avalon_sdcard_slave_read;                                    // mm_interconnect_0:SD_Card_avalon_sdcard_slave_read -> SD_Card:i_avalon_read
	wire   [3:0] mm_interconnect_0_sd_card_avalon_sdcard_slave_byteenable;                              // mm_interconnect_0:SD_Card_avalon_sdcard_slave_byteenable -> SD_Card:i_avalon_byteenable
	wire         mm_interconnect_0_sd_card_avalon_sdcard_slave_write;                                   // mm_interconnect_0:SD_Card_avalon_sdcard_slave_write -> SD_Card:i_avalon_write
	wire  [31:0] mm_interconnect_0_sd_card_avalon_sdcard_slave_writedata;                               // mm_interconnect_0:SD_Card_avalon_sdcard_slave_writedata -> SD_Card:i_avalon_writedata
	wire  [15:0] mm_interconnect_0_sram_avalon_sram_slave_readdata;                                     // SRAM:readdata -> mm_interconnect_0:SRAM_avalon_sram_slave_readdata
	wire  [19:0] mm_interconnect_0_sram_avalon_sram_slave_address;                                      // mm_interconnect_0:SRAM_avalon_sram_slave_address -> SRAM:address
	wire         mm_interconnect_0_sram_avalon_sram_slave_read;                                         // mm_interconnect_0:SRAM_avalon_sram_slave_read -> SRAM:read
	wire   [1:0] mm_interconnect_0_sram_avalon_sram_slave_byteenable;                                   // mm_interconnect_0:SRAM_avalon_sram_slave_byteenable -> SRAM:byteenable
	wire         mm_interconnect_0_sram_avalon_sram_slave_readdatavalid;                                // SRAM:readdatavalid -> mm_interconnect_0:SRAM_avalon_sram_slave_readdatavalid
	wire         mm_interconnect_0_sram_avalon_sram_slave_write;                                        // mm_interconnect_0:SRAM_avalon_sram_slave_write -> SRAM:write
	wire  [15:0] mm_interconnect_0_sram_avalon_sram_slave_writedata;                                    // mm_interconnect_0:SRAM_avalon_sram_slave_writedata -> SRAM:writedata
	wire         mm_interconnect_0_usb_avalon_usb_slave_chipselect;                                     // mm_interconnect_0:USB_avalon_usb_slave_chipselect -> USB:chipselect
	wire  [15:0] mm_interconnect_0_usb_avalon_usb_slave_readdata;                                       // USB:readdata -> mm_interconnect_0:USB_avalon_usb_slave_readdata
	wire   [1:0] mm_interconnect_0_usb_avalon_usb_slave_address;                                        // mm_interconnect_0:USB_avalon_usb_slave_address -> USB:address
	wire         mm_interconnect_0_usb_avalon_usb_slave_read;                                           // mm_interconnect_0:USB_avalon_usb_slave_read -> USB:read
	wire         mm_interconnect_0_usb_avalon_usb_slave_write;                                          // mm_interconnect_0:USB_avalon_usb_slave_write -> USB:write
	wire  [15:0] mm_interconnect_0_usb_avalon_usb_slave_writedata;                                      // mm_interconnect_0:USB_avalon_usb_slave_writedata -> USB:writedata
	wire  [31:0] mm_interconnect_0_vga_subsystem_char_buffer_control_slave_readdata;                    // VGA_Subsystem:char_buffer_control_slave_readdata -> mm_interconnect_0:VGA_Subsystem_char_buffer_control_slave_readdata
	wire   [1:0] mm_interconnect_0_vga_subsystem_char_buffer_control_slave_address;                     // mm_interconnect_0:VGA_Subsystem_char_buffer_control_slave_address -> VGA_Subsystem:char_buffer_control_slave_address
	wire         mm_interconnect_0_vga_subsystem_char_buffer_control_slave_read;                        // mm_interconnect_0:VGA_Subsystem_char_buffer_control_slave_read -> VGA_Subsystem:char_buffer_control_slave_read
	wire   [3:0] mm_interconnect_0_vga_subsystem_char_buffer_control_slave_byteenable;                  // mm_interconnect_0:VGA_Subsystem_char_buffer_control_slave_byteenable -> VGA_Subsystem:char_buffer_control_slave_byteenable
	wire         mm_interconnect_0_vga_subsystem_char_buffer_control_slave_write;                       // mm_interconnect_0:VGA_Subsystem_char_buffer_control_slave_write -> VGA_Subsystem:char_buffer_control_slave_write
	wire  [31:0] mm_interconnect_0_vga_subsystem_char_buffer_control_slave_writedata;                   // mm_interconnect_0:VGA_Subsystem_char_buffer_control_slave_writedata -> VGA_Subsystem:char_buffer_control_slave_writedata
	wire         mm_interconnect_0_vga_subsystem_char_buffer_slave_chipselect;                          // mm_interconnect_0:VGA_Subsystem_char_buffer_slave_chipselect -> VGA_Subsystem:char_buffer_slave_chipselect
	wire  [31:0] mm_interconnect_0_vga_subsystem_char_buffer_slave_readdata;                            // VGA_Subsystem:char_buffer_slave_readdata -> mm_interconnect_0:VGA_Subsystem_char_buffer_slave_readdata
	wire  [10:0] mm_interconnect_0_vga_subsystem_char_buffer_slave_address;                             // mm_interconnect_0:VGA_Subsystem_char_buffer_slave_address -> VGA_Subsystem:char_buffer_slave_address
	wire   [3:0] mm_interconnect_0_vga_subsystem_char_buffer_slave_byteenable;                          // mm_interconnect_0:VGA_Subsystem_char_buffer_slave_byteenable -> VGA_Subsystem:char_buffer_slave_byteenable
	wire         mm_interconnect_0_vga_subsystem_char_buffer_slave_write;                               // mm_interconnect_0:VGA_Subsystem_char_buffer_slave_write -> VGA_Subsystem:char_buffer_slave_write
	wire  [31:0] mm_interconnect_0_vga_subsystem_char_buffer_slave_writedata;                           // mm_interconnect_0:VGA_Subsystem_char_buffer_slave_writedata -> VGA_Subsystem:char_buffer_slave_writedata
	wire         mm_interconnect_0_vga_subsystem_char_buffer_slave_clken;                               // mm_interconnect_0:VGA_Subsystem_char_buffer_slave_clken -> VGA_Subsystem:char_buffer_slave_clken
	wire  [31:0] mm_interconnect_0_sysid_control_slave_readdata;                                        // SysID:readdata -> mm_interconnect_0:SysID_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_control_slave_address;                                         // mm_interconnect_0:SysID_control_slave_address -> SysID:address
	wire  [31:0] mm_interconnect_0_nios2_debug_mem_slave_readdata;                                      // Nios2:debug_mem_slave_readdata -> mm_interconnect_0:Nios2_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_debug_mem_slave_waitrequest;                                   // Nios2:debug_mem_slave_waitrequest -> mm_interconnect_0:Nios2_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_debug_mem_slave_debugaccess;                                   // mm_interconnect_0:Nios2_debug_mem_slave_debugaccess -> Nios2:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_debug_mem_slave_address;                                       // mm_interconnect_0:Nios2_debug_mem_slave_address -> Nios2:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_debug_mem_slave_read;                                          // mm_interconnect_0:Nios2_debug_mem_slave_read -> Nios2:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_debug_mem_slave_byteenable;                                    // mm_interconnect_0:Nios2_debug_mem_slave_byteenable -> Nios2:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_debug_mem_slave_write;                                         // mm_interconnect_0:Nios2_debug_mem_slave_write -> Nios2:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_debug_mem_slave_writedata;                                     // mm_interconnect_0:Nios2_debug_mem_slave_writedata -> Nios2:debug_mem_slave_writedata
	wire         mm_interconnect_0_flash_flash_data_chipselect;                                         // mm_interconnect_0:Flash_flash_data_chipselect -> Flash:i_avalon_chip_select
	wire  [31:0] mm_interconnect_0_flash_flash_data_readdata;                                           // Flash:o_avalon_readdata -> mm_interconnect_0:Flash_flash_data_readdata
	wire         mm_interconnect_0_flash_flash_data_waitrequest;                                        // Flash:o_avalon_waitrequest -> mm_interconnect_0:Flash_flash_data_waitrequest
	wire  [20:0] mm_interconnect_0_flash_flash_data_address;                                            // mm_interconnect_0:Flash_flash_data_address -> Flash:i_avalon_address
	wire         mm_interconnect_0_flash_flash_data_read;                                               // mm_interconnect_0:Flash_flash_data_read -> Flash:i_avalon_read
	wire   [3:0] mm_interconnect_0_flash_flash_data_byteenable;                                         // mm_interconnect_0:Flash_flash_data_byteenable -> Flash:i_avalon_byteenable
	wire         mm_interconnect_0_flash_flash_data_write;                                              // mm_interconnect_0:Flash_flash_data_write -> Flash:i_avalon_write
	wire  [31:0] mm_interconnect_0_flash_flash_data_writedata;                                          // mm_interconnect_0:Flash_flash_data_writedata -> Flash:i_avalon_writedata
	wire         mm_interconnect_0_flash_flash_erase_control_chipselect;                                // mm_interconnect_0:Flash_flash_erase_control_chipselect -> Flash:i_avalon_erase_chip_select
	wire  [31:0] mm_interconnect_0_flash_flash_erase_control_readdata;                                  // Flash:o_avalon_erase_readdata -> mm_interconnect_0:Flash_flash_erase_control_readdata
	wire         mm_interconnect_0_flash_flash_erase_control_waitrequest;                               // Flash:o_avalon_erase_waitrequest -> mm_interconnect_0:Flash_flash_erase_control_waitrequest
	wire         mm_interconnect_0_flash_flash_erase_control_read;                                      // mm_interconnect_0:Flash_flash_erase_control_read -> Flash:i_avalon_erase_read
	wire   [3:0] mm_interconnect_0_flash_flash_erase_control_byteenable;                                // mm_interconnect_0:Flash_flash_erase_control_byteenable -> Flash:i_avalon_erase_byteenable
	wire         mm_interconnect_0_flash_flash_erase_control_write;                                     // mm_interconnect_0:Flash_flash_erase_control_write -> Flash:i_avalon_erase_write
	wire  [31:0] mm_interconnect_0_flash_flash_erase_control_writedata;                                 // mm_interconnect_0:Flash_flash_erase_control_writedata -> Flash:i_avalon_erase_writedata
	wire  [31:0] mm_interconnect_0_vga_subsystem_pixel_dma_control_slave_readdata;                      // VGA_Subsystem:pixel_dma_control_slave_readdata -> mm_interconnect_0:VGA_Subsystem_pixel_dma_control_slave_readdata
	wire   [1:0] mm_interconnect_0_vga_subsystem_pixel_dma_control_slave_address;                       // mm_interconnect_0:VGA_Subsystem_pixel_dma_control_slave_address -> VGA_Subsystem:pixel_dma_control_slave_address
	wire         mm_interconnect_0_vga_subsystem_pixel_dma_control_slave_read;                          // mm_interconnect_0:VGA_Subsystem_pixel_dma_control_slave_read -> VGA_Subsystem:pixel_dma_control_slave_read
	wire   [3:0] mm_interconnect_0_vga_subsystem_pixel_dma_control_slave_byteenable;                    // mm_interconnect_0:VGA_Subsystem_pixel_dma_control_slave_byteenable -> VGA_Subsystem:pixel_dma_control_slave_byteenable
	wire         mm_interconnect_0_vga_subsystem_pixel_dma_control_slave_write;                         // mm_interconnect_0:VGA_Subsystem_pixel_dma_control_slave_write -> VGA_Subsystem:pixel_dma_control_slave_write
	wire  [31:0] mm_interconnect_0_vga_subsystem_pixel_dma_control_slave_writedata;                     // mm_interconnect_0:VGA_Subsystem_pixel_dma_control_slave_writedata -> VGA_Subsystem:pixel_dma_control_slave_writedata
	wire  [31:0] mm_interconnect_0_vga_subsystem_rgb_slave_readdata;                                    // VGA_Subsystem:rgb_slave_readdata -> mm_interconnect_0:VGA_Subsystem_rgb_slave_readdata
	wire         mm_interconnect_0_vga_subsystem_rgb_slave_read;                                        // mm_interconnect_0:VGA_Subsystem_rgb_slave_read -> VGA_Subsystem:rgb_slave_read
	wire         mm_interconnect_0_sdram_s1_chipselect;                                                 // mm_interconnect_0:SDRAM_s1_chipselect -> SDRAM:az_cs
	wire  [31:0] mm_interconnect_0_sdram_s1_readdata;                                                   // SDRAM:za_data -> mm_interconnect_0:SDRAM_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;                                                // SDRAM:za_waitrequest -> mm_interconnect_0:SDRAM_s1_waitrequest
	wire  [24:0] mm_interconnect_0_sdram_s1_address;                                                    // mm_interconnect_0:SDRAM_s1_address -> SDRAM:az_addr
	wire         mm_interconnect_0_sdram_s1_read;                                                       // mm_interconnect_0:SDRAM_s1_read -> SDRAM:az_rd_n
	wire   [3:0] mm_interconnect_0_sdram_s1_byteenable;                                                 // mm_interconnect_0:SDRAM_s1_byteenable -> SDRAM:az_be_n
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                                              // SDRAM:za_valid -> mm_interconnect_0:SDRAM_s1_readdatavalid
	wire         mm_interconnect_0_sdram_s1_write;                                                      // mm_interconnect_0:SDRAM_s1_write -> SDRAM:az_wr_n
	wire  [31:0] mm_interconnect_0_sdram_s1_writedata;                                                  // mm_interconnect_0:SDRAM_s1_writedata -> SDRAM:az_data
	wire         mm_interconnect_0_red_leds_s1_chipselect;                                              // mm_interconnect_0:Red_LEDs_s1_chipselect -> Red_LEDs:chipselect
	wire  [31:0] mm_interconnect_0_red_leds_s1_readdata;                                                // Red_LEDs:readdata -> mm_interconnect_0:Red_LEDs_s1_readdata
	wire   [1:0] mm_interconnect_0_red_leds_s1_address;                                                 // mm_interconnect_0:Red_LEDs_s1_address -> Red_LEDs:address
	wire         mm_interconnect_0_red_leds_s1_write;                                                   // mm_interconnect_0:Red_LEDs_s1_write -> Red_LEDs:write_n
	wire  [31:0] mm_interconnect_0_red_leds_s1_writedata;                                               // mm_interconnect_0:Red_LEDs_s1_writedata -> Red_LEDs:writedata
	wire         mm_interconnect_0_green_leds_s1_chipselect;                                            // mm_interconnect_0:Green_LEDs_s1_chipselect -> Green_LEDs:chipselect
	wire  [31:0] mm_interconnect_0_green_leds_s1_readdata;                                              // Green_LEDs:readdata -> mm_interconnect_0:Green_LEDs_s1_readdata
	wire   [1:0] mm_interconnect_0_green_leds_s1_address;                                               // mm_interconnect_0:Green_LEDs_s1_address -> Green_LEDs:address
	wire         mm_interconnect_0_green_leds_s1_write;                                                 // mm_interconnect_0:Green_LEDs_s1_write -> Green_LEDs:write_n
	wire  [31:0] mm_interconnect_0_green_leds_s1_writedata;                                             // mm_interconnect_0:Green_LEDs_s1_writedata -> Green_LEDs:writedata
	wire         mm_interconnect_0_hex3_hex0_s1_chipselect;                                             // mm_interconnect_0:HEX3_HEX0_s1_chipselect -> HEX3_HEX0:chipselect
	wire  [31:0] mm_interconnect_0_hex3_hex0_s1_readdata;                                               // HEX3_HEX0:readdata -> mm_interconnect_0:HEX3_HEX0_s1_readdata
	wire   [1:0] mm_interconnect_0_hex3_hex0_s1_address;                                                // mm_interconnect_0:HEX3_HEX0_s1_address -> HEX3_HEX0:address
	wire         mm_interconnect_0_hex3_hex0_s1_write;                                                  // mm_interconnect_0:HEX3_HEX0_s1_write -> HEX3_HEX0:write_n
	wire  [31:0] mm_interconnect_0_hex3_hex0_s1_writedata;                                              // mm_interconnect_0:HEX3_HEX0_s1_writedata -> HEX3_HEX0:writedata
	wire         mm_interconnect_0_hex7_hex4_s1_chipselect;                                             // mm_interconnect_0:HEX7_HEX4_s1_chipselect -> HEX7_HEX4:chipselect
	wire  [31:0] mm_interconnect_0_hex7_hex4_s1_readdata;                                               // HEX7_HEX4:readdata -> mm_interconnect_0:HEX7_HEX4_s1_readdata
	wire   [1:0] mm_interconnect_0_hex7_hex4_s1_address;                                                // mm_interconnect_0:HEX7_HEX4_s1_address -> HEX7_HEX4:address
	wire         mm_interconnect_0_hex7_hex4_s1_write;                                                  // mm_interconnect_0:HEX7_HEX4_s1_write -> HEX7_HEX4:write_n
	wire  [31:0] mm_interconnect_0_hex7_hex4_s1_writedata;                                              // mm_interconnect_0:HEX7_HEX4_s1_writedata -> HEX7_HEX4:writedata
	wire  [31:0] mm_interconnect_0_slider_switches_s1_readdata;                                         // Slider_Switches:readdata -> mm_interconnect_0:Slider_Switches_s1_readdata
	wire   [1:0] mm_interconnect_0_slider_switches_s1_address;                                          // mm_interconnect_0:Slider_Switches_s1_address -> Slider_Switches:address
	wire         mm_interconnect_0_pushbuttons_s1_chipselect;                                           // mm_interconnect_0:Pushbuttons_s1_chipselect -> Pushbuttons:chipselect
	wire  [31:0] mm_interconnect_0_pushbuttons_s1_readdata;                                             // Pushbuttons:readdata -> mm_interconnect_0:Pushbuttons_s1_readdata
	wire   [1:0] mm_interconnect_0_pushbuttons_s1_address;                                              // mm_interconnect_0:Pushbuttons_s1_address -> Pushbuttons:address
	wire         mm_interconnect_0_pushbuttons_s1_write;                                                // mm_interconnect_0:Pushbuttons_s1_write -> Pushbuttons:write_n
	wire  [31:0] mm_interconnect_0_pushbuttons_s1_writedata;                                            // mm_interconnect_0:Pushbuttons_s1_writedata -> Pushbuttons:writedata
	wire         mm_interconnect_0_expansion_jp5_s1_chipselect;                                         // mm_interconnect_0:Expansion_JP5_s1_chipselect -> Expansion_JP5:chipselect
	wire  [31:0] mm_interconnect_0_expansion_jp5_s1_readdata;                                           // Expansion_JP5:readdata -> mm_interconnect_0:Expansion_JP5_s1_readdata
	wire   [1:0] mm_interconnect_0_expansion_jp5_s1_address;                                            // mm_interconnect_0:Expansion_JP5_s1_address -> Expansion_JP5:address
	wire         mm_interconnect_0_expansion_jp5_s1_write;                                              // mm_interconnect_0:Expansion_JP5_s1_write -> Expansion_JP5:write_n
	wire  [31:0] mm_interconnect_0_expansion_jp5_s1_writedata;                                          // mm_interconnect_0:Expansion_JP5_s1_writedata -> Expansion_JP5:writedata
	wire         mm_interconnect_0_interval_timer_s1_chipselect;                                        // mm_interconnect_0:Interval_Timer_s1_chipselect -> Interval_Timer:chipselect
	wire  [15:0] mm_interconnect_0_interval_timer_s1_readdata;                                          // Interval_Timer:readdata -> mm_interconnect_0:Interval_Timer_s1_readdata
	wire   [2:0] mm_interconnect_0_interval_timer_s1_address;                                           // mm_interconnect_0:Interval_Timer_s1_address -> Interval_Timer:address
	wire         mm_interconnect_0_interval_timer_s1_write;                                             // mm_interconnect_0:Interval_Timer_s1_write -> Interval_Timer:write_n
	wire  [15:0] mm_interconnect_0_interval_timer_s1_writedata;                                         // mm_interconnect_0:Interval_Timer_s1_writedata -> Interval_Timer:writedata
	wire         mm_interconnect_0_interval_timer_2_s1_chipselect;                                      // mm_interconnect_0:Interval_Timer_2_s1_chipselect -> Interval_Timer_2:chipselect
	wire  [15:0] mm_interconnect_0_interval_timer_2_s1_readdata;                                        // Interval_Timer_2:readdata -> mm_interconnect_0:Interval_Timer_2_s1_readdata
	wire   [2:0] mm_interconnect_0_interval_timer_2_s1_address;                                         // mm_interconnect_0:Interval_Timer_2_s1_address -> Interval_Timer_2:address
	wire         mm_interconnect_0_interval_timer_2_s1_write;                                           // mm_interconnect_0:Interval_Timer_2_s1_write -> Interval_Timer_2:write_n
	wire  [15:0] mm_interconnect_0_interval_timer_2_s1_writedata;                                       // mm_interconnect_0:Interval_Timer_2_s1_writedata -> Interval_Timer_2:writedata
	wire  [31:0] mm_interconnect_0_video_in_subsystem_video_in_dma_control_slave_readdata;              // Video_In_Subsystem:video_in_dma_control_slave_readdata -> mm_interconnect_0:Video_In_Subsystem_video_in_dma_control_slave_readdata
	wire   [1:0] mm_interconnect_0_video_in_subsystem_video_in_dma_control_slave_address;               // mm_interconnect_0:Video_In_Subsystem_video_in_dma_control_slave_address -> Video_In_Subsystem:video_in_dma_control_slave_address
	wire         mm_interconnect_0_video_in_subsystem_video_in_dma_control_slave_read;                  // mm_interconnect_0:Video_In_Subsystem_video_in_dma_control_slave_read -> Video_In_Subsystem:video_in_dma_control_slave_read
	wire   [3:0] mm_interconnect_0_video_in_subsystem_video_in_dma_control_slave_byteenable;            // mm_interconnect_0:Video_In_Subsystem_video_in_dma_control_slave_byteenable -> Video_In_Subsystem:video_in_dma_control_slave_byteenable
	wire         mm_interconnect_0_video_in_subsystem_video_in_dma_control_slave_write;                 // mm_interconnect_0:Video_In_Subsystem_video_in_dma_control_slave_write -> Video_In_Subsystem:video_in_dma_control_slave_write
	wire  [31:0] mm_interconnect_0_video_in_subsystem_video_in_dma_control_slave_writedata;             // mm_interconnect_0:Video_In_Subsystem_video_in_dma_control_slave_writedata -> Video_In_Subsystem:video_in_dma_control_slave_writedata
	wire         mm_interconnect_0_video_in_subsystem_video_in_edge_detection_control_slave_chipselect; // mm_interconnect_0:Video_In_Subsystem_video_in_edge_detection_control_slave_chipselect -> Video_In_Subsystem:video_in_edge_detection_control_slave_chipselect
	wire  [31:0] mm_interconnect_0_video_in_subsystem_video_in_edge_detection_control_slave_readdata;   // Video_In_Subsystem:video_in_edge_detection_control_slave_readdata -> mm_interconnect_0:Video_In_Subsystem_video_in_edge_detection_control_slave_readdata
	wire   [1:0] mm_interconnect_0_video_in_subsystem_video_in_edge_detection_control_slave_address;    // mm_interconnect_0:Video_In_Subsystem_video_in_edge_detection_control_slave_address -> Video_In_Subsystem:video_in_edge_detection_control_slave_address
	wire         mm_interconnect_0_video_in_subsystem_video_in_edge_detection_control_slave_write;      // mm_interconnect_0:Video_In_Subsystem_video_in_edge_detection_control_slave_write -> Video_In_Subsystem:video_in_edge_detection_control_slave_write_n
	wire  [31:0] mm_interconnect_0_video_in_subsystem_video_in_edge_detection_control_slave_writedata;  // mm_interconnect_0:Video_In_Subsystem_video_in_edge_detection_control_slave_writedata -> Video_In_Subsystem:video_in_edge_detection_control_slave_writedata
	wire         mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_chipselect;                     // mm_interconnect_0:JTAG_UART_2nd_Core_avalon_jtag_slave_chipselect -> JTAG_UART_2nd_Core:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_readdata;                       // JTAG_UART_2nd_Core:av_readdata -> mm_interconnect_0:JTAG_UART_2nd_Core_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_waitrequest;                    // JTAG_UART_2nd_Core:av_waitrequest -> mm_interconnect_0:JTAG_UART_2nd_Core_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_address;                        // mm_interconnect_0:JTAG_UART_2nd_Core_avalon_jtag_slave_address -> JTAG_UART_2nd_Core:av_address
	wire         mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_read;                           // mm_interconnect_0:JTAG_UART_2nd_Core_avalon_jtag_slave_read -> JTAG_UART_2nd_Core:av_read_n
	wire         mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_write;                          // mm_interconnect_0:JTAG_UART_2nd_Core_avalon_jtag_slave_write -> JTAG_UART_2nd_Core:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_writedata;                      // mm_interconnect_0:JTAG_UART_2nd_Core_avalon_jtag_slave_writedata -> JTAG_UART_2nd_Core:av_writedata
	wire  [31:0] mm_interconnect_0_nios2_2nd_core_debug_mem_slave_readdata;                             // Nios2_2nd_Core:debug_mem_slave_readdata -> mm_interconnect_0:Nios2_2nd_Core_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_2nd_core_debug_mem_slave_waitrequest;                          // Nios2_2nd_Core:debug_mem_slave_waitrequest -> mm_interconnect_0:Nios2_2nd_Core_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_2nd_core_debug_mem_slave_debugaccess;                          // mm_interconnect_0:Nios2_2nd_Core_debug_mem_slave_debugaccess -> Nios2_2nd_Core:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_2nd_core_debug_mem_slave_address;                              // mm_interconnect_0:Nios2_2nd_Core_debug_mem_slave_address -> Nios2_2nd_Core:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_2nd_core_debug_mem_slave_read;                                 // mm_interconnect_0:Nios2_2nd_Core_debug_mem_slave_read -> Nios2_2nd_Core:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_2nd_core_debug_mem_slave_byteenable;                           // mm_interconnect_0:Nios2_2nd_Core_debug_mem_slave_byteenable -> Nios2_2nd_Core:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_2nd_core_debug_mem_slave_write;                                // mm_interconnect_0:Nios2_2nd_Core_debug_mem_slave_write -> Nios2_2nd_Core:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_2nd_core_debug_mem_slave_writedata;                            // mm_interconnect_0:Nios2_2nd_Core_debug_mem_slave_writedata -> Nios2_2nd_Core:debug_mem_slave_writedata
	wire         mm_interconnect_0_interval_timer_2nd_core_s1_chipselect;                               // mm_interconnect_0:Interval_Timer_2nd_Core_s1_chipselect -> Interval_Timer_2nd_Core:chipselect
	wire  [15:0] mm_interconnect_0_interval_timer_2nd_core_s1_readdata;                                 // Interval_Timer_2nd_Core:readdata -> mm_interconnect_0:Interval_Timer_2nd_Core_s1_readdata
	wire   [2:0] mm_interconnect_0_interval_timer_2nd_core_s1_address;                                  // mm_interconnect_0:Interval_Timer_2nd_Core_s1_address -> Interval_Timer_2nd_Core:address
	wire         mm_interconnect_0_interval_timer_2nd_core_s1_write;                                    // mm_interconnect_0:Interval_Timer_2nd_Core_s1_write -> Interval_Timer_2nd_Core:write_n
	wire  [15:0] mm_interconnect_0_interval_timer_2nd_core_s1_writedata;                                // mm_interconnect_0:Interval_Timer_2nd_Core_s1_writedata -> Interval_Timer_2nd_Core:writedata
	wire         mm_interconnect_0_interval_timer_2nd_core_2_s1_chipselect;                             // mm_interconnect_0:Interval_Timer_2nd_Core_2_s1_chipselect -> Interval_Timer_2nd_Core_2:chipselect
	wire  [15:0] mm_interconnect_0_interval_timer_2nd_core_2_s1_readdata;                               // Interval_Timer_2nd_Core_2:readdata -> mm_interconnect_0:Interval_Timer_2nd_Core_2_s1_readdata
	wire   [2:0] mm_interconnect_0_interval_timer_2nd_core_2_s1_address;                                // mm_interconnect_0:Interval_Timer_2nd_Core_2_s1_address -> Interval_Timer_2nd_Core_2:address
	wire         mm_interconnect_0_interval_timer_2nd_core_2_s1_write;                                  // mm_interconnect_0:Interval_Timer_2nd_Core_2_s1_write -> Interval_Timer_2nd_Core_2:write_n
	wire  [15:0] mm_interconnect_0_interval_timer_2nd_core_2_s1_writedata;                              // mm_interconnect_0:Interval_Timer_2nd_Core_2_s1_writedata -> Interval_Timer_2nd_Core_2:writedata
	wire         irq_mapper_receiver8_irq;                                                              // JTAG_UART:av_irq -> irq_mapper:receiver8_irq
	wire         irq_mapper_receiver9_irq;                                                              // Interval_Timer:irq -> irq_mapper:receiver9_irq
	wire         irq_mapper_receiver10_irq;                                                             // Interval_Timer_2:irq -> irq_mapper:receiver10_irq
	wire  [31:0] nios2_irq_irq;                                                                         // irq_mapper:sender_irq -> Nios2:irq
	wire         irq_mapper_001_receiver8_irq;                                                          // JTAG_UART_2nd_Core:av_irq -> irq_mapper_001:receiver8_irq
	wire         irq_mapper_001_receiver9_irq;                                                          // Interval_Timer_2nd_Core:irq -> irq_mapper_001:receiver9_irq
	wire         irq_mapper_001_receiver10_irq;                                                         // Interval_Timer_2nd_Core_2:irq -> irq_mapper_001:receiver10_irq
	wire  [31:0] nios2_2nd_core_irq_irq;                                                                // irq_mapper_001:sender_irq -> Nios2_2nd_Core:irq
	wire         irq_mapper_receiver0_irq;                                                              // Audio_Subsystem:audio_irq_irq -> [irq_mapper:receiver0_irq, irq_mapper_001:receiver0_irq]
	wire         irq_mapper_receiver7_irq;                                                              // Expansion_JP5:irq -> [irq_mapper:receiver7_irq, irq_mapper_001:receiver7_irq]
	wire         irq_mapper_receiver5_irq;                                                              // IrDA:irq -> [irq_mapper:receiver5_irq, irq_mapper_001:receiver5_irq]
	wire         irq_mapper_receiver1_irq;                                                              // PS2_Port:irq -> [irq_mapper:receiver1_irq, irq_mapper_001:receiver1_irq]
	wire         irq_mapper_receiver2_irq;                                                              // PS2_Port_Dual:irq -> [irq_mapper:receiver2_irq, irq_mapper_001:receiver2_irq]
	wire         irq_mapper_receiver6_irq;                                                              // Pushbuttons:irq -> [irq_mapper:receiver6_irq, irq_mapper_001:receiver6_irq]
	wire         irq_mapper_receiver4_irq;                                                              // Serial_Port:irq -> [irq_mapper:receiver4_irq, irq_mapper_001:receiver4_irq]
	wire         irq_mapper_receiver3_irq;                                                              // USB:irq -> [irq_mapper:receiver3_irq, irq_mapper_001:receiver3_irq]
	wire         rst_controller_reset_out_reset;                                                        // rst_controller:reset_out -> [AV_Config:reset, Char_LCD_16x2:reset, Expansion_JP5:reset_n, Flash:i_reset_n, Green_LEDs:reset_n, HEX3_HEX0:reset_n, HEX7_HEX4:reset_n, Interval_Timer:reset_n, Interval_Timer_2:reset_n, Interval_Timer_2nd_Core:reset_n, Interval_Timer_2nd_Core_2:reset_n, IrDA:reset, JTAG_UART:rst_n, JTAG_UART_2nd_Core:rst_n, PS2_Port:reset, PS2_Port_Dual:reset, Pushbuttons:reset_n, Red_LEDs:reset_n, SDRAM:reset_n, SD_Card:i_reset_n, SRAM:reset, Serial_Port:reset, Slider_Switches:reset_n, SysID:reset_n, USB:reset, mm_interconnect_0:AV_Config_reset_reset_bridge_in_reset_reset, mm_interconnect_0:JTAG_to_FPGA_Bridge_clk_reset_reset_bridge_in_reset_reset]
	wire         rst_controller_001_reset_out_reset;                                                    // rst_controller_001:reset_out -> [Nios2:reset_n, irq_mapper:reset, mm_interconnect_0:Nios2_reset_reset_bridge_in_reset_reset]
	wire         nios2_debug_reset_request_reset;                                                       // Nios2:debug_reset_request -> rst_controller_001:reset_in0
	wire         rst_controller_002_reset_out_reset;                                                    // rst_controller_002:reset_out -> [Nios2_2nd_Core:reset_n, irq_mapper_001:reset, mm_interconnect_0:Nios2_2nd_Core_reset_reset_bridge_in_reset_reset]
	wire         nios2_2nd_core_debug_reset_request_reset;                                              // Nios2_2nd_Core:debug_reset_request -> rst_controller_002:reset_in0

	Computer_System_AV_Config av_config (
		.clk         (system_pll_sys_clk_clk),                                         //                    clk.clk
		.reset       (rst_controller_reset_out_reset),                                 //                  reset.reset
		.address     (mm_interconnect_0_av_config_avalon_av_config_slave_address),     // avalon_av_config_slave.address
		.byteenable  (mm_interconnect_0_av_config_avalon_av_config_slave_byteenable),  //                       .byteenable
		.read        (mm_interconnect_0_av_config_avalon_av_config_slave_read),        //                       .read
		.write       (mm_interconnect_0_av_config_avalon_av_config_slave_write),       //                       .write
		.writedata   (mm_interconnect_0_av_config_avalon_av_config_slave_writedata),   //                       .writedata
		.readdata    (mm_interconnect_0_av_config_avalon_av_config_slave_readdata),    //                       .readdata
		.waitrequest (mm_interconnect_0_av_config_avalon_av_config_slave_waitrequest), //                       .waitrequest
		.I2C_SDAT    (av_config_SDAT),                                                 //     external_interface.export
		.I2C_SCLK    (av_config_SCLK)                                                  //                       .export
	);

	Computer_System_Audio_Subsystem audio_subsystem (
		.audio_ADCDAT              (audio_ADCDAT),                                             //               audio.ADCDAT
		.audio_ADCLRCK             (audio_ADCLRCK),                                            //                    .ADCLRCK
		.audio_BCLK                (audio_BCLK),                                               //                    .BCLK
		.audio_DACDAT              (audio_DACDAT),                                             //                    .DACDAT
		.audio_DACLRCK             (audio_DACLRCK),                                            //                    .DACLRCK
		.audio_irq_irq             (irq_mapper_receiver0_irq),                                 //           audio_irq.irq
		.audio_pll_clk_clk         (audio_pll_clk_clk),                                        //       audio_pll_clk.clk
		.audio_pll_ref_clk_clk     (audio_pll_ref_clk_clk),                                    //   audio_pll_ref_clk.clk
		.audio_pll_ref_reset_reset (audio_pll_ref_reset_reset),                                // audio_pll_ref_reset.reset
		.audio_pll_reset_reset     (),                                                         //     audio_pll_reset.reset
		.audio_slave_address       (mm_interconnect_0_audio_subsystem_audio_slave_address),    //         audio_slave.address
		.audio_slave_chipselect    (mm_interconnect_0_audio_subsystem_audio_slave_chipselect), //                    .chipselect
		.audio_slave_read          (mm_interconnect_0_audio_subsystem_audio_slave_read),       //                    .read
		.audio_slave_write         (mm_interconnect_0_audio_subsystem_audio_slave_write),      //                    .write
		.audio_slave_writedata     (mm_interconnect_0_audio_subsystem_audio_slave_writedata),  //                    .writedata
		.audio_slave_readdata      (mm_interconnect_0_audio_subsystem_audio_slave_readdata),   //                    .readdata
		.sys_clk_clk               (system_pll_sys_clk_clk),                                   //             sys_clk.clk
		.sys_reset_reset_n         (~system_pll_reset_source_reset)                            //           sys_reset.reset_n
	);

	Computer_System_Char_LCD_16x2 char_lcd_16x2 (
		.clk         (system_pll_sys_clk_clk),                                       //                clk.clk
		.reset       (rst_controller_reset_out_reset),                               //              reset.reset
		.address     (mm_interconnect_0_char_lcd_16x2_avalon_lcd_slave_address),     //   avalon_lcd_slave.address
		.chipselect  (mm_interconnect_0_char_lcd_16x2_avalon_lcd_slave_chipselect),  //                   .chipselect
		.read        (mm_interconnect_0_char_lcd_16x2_avalon_lcd_slave_read),        //                   .read
		.write       (mm_interconnect_0_char_lcd_16x2_avalon_lcd_slave_write),       //                   .write
		.writedata   (mm_interconnect_0_char_lcd_16x2_avalon_lcd_slave_writedata),   //                   .writedata
		.readdata    (mm_interconnect_0_char_lcd_16x2_avalon_lcd_slave_readdata),    //                   .readdata
		.waitrequest (mm_interconnect_0_char_lcd_16x2_avalon_lcd_slave_waitrequest), //                   .waitrequest
		.LCD_DATA    (char_lcd_DATA),                                                // external_interface.export
		.LCD_ON      (char_lcd_ON),                                                  //                   .export
		.LCD_BLON    (char_lcd_BLON),                                                //                   .export
		.LCD_EN      (char_lcd_EN),                                                  //                   .export
		.LCD_RS      (char_lcd_RS),                                                  //                   .export
		.LCD_RW      (char_lcd_RW)                                                   //                   .export
	);

	Computer_System_Expansion_JP5 expansion_jp5 (
		.clk        (system_pll_sys_clk_clk),                        //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address    (mm_interconnect_0_expansion_jp5_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_expansion_jp5_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_expansion_jp5_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_expansion_jp5_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_expansion_jp5_s1_readdata),   //                    .readdata
		.bidir_port (expansion_jp5_export),                          // external_connection.export
		.irq        (irq_mapper_receiver7_irq)                       //                 irq.irq
	);

	Altera_UP_Flash_Memory_IP_Core_Avalon_Interface #(
		.FLASH_MEMORY_ADDRESS_WIDTH (23)
	) flash (
		.i_avalon_chip_select       (mm_interconnect_0_flash_flash_data_chipselect),           //          flash_data.chipselect
		.i_avalon_write             (mm_interconnect_0_flash_flash_data_write),                //                    .write
		.i_avalon_read              (mm_interconnect_0_flash_flash_data_read),                 //                    .read
		.i_avalon_address           (mm_interconnect_0_flash_flash_data_address),              //                    .address
		.i_avalon_byteenable        (mm_interconnect_0_flash_flash_data_byteenable),           //                    .byteenable
		.i_avalon_writedata         (mm_interconnect_0_flash_flash_data_writedata),            //                    .writedata
		.o_avalon_readdata          (mm_interconnect_0_flash_flash_data_readdata),             //                    .readdata
		.o_avalon_waitrequest       (mm_interconnect_0_flash_flash_data_waitrequest),          //                    .waitrequest
		.i_clock                    (system_pll_sys_clk_clk),                                  //                 clk.clk
		.i_reset_n                  (~rst_controller_reset_out_reset),                         //               reset.reset_n
		.FL_ADDR                    (flash_ADDR),                                              //         conduit_end.export
		.FL_CE_N                    (flash_CE_N),                                              //                    .export
		.FL_OE_N                    (flash_OE_N),                                              //                    .export
		.FL_WE_N                    (flash_WE_N),                                              //                    .export
		.FL_RST_N                   (flash_RST_N),                                             //                    .export
		.FL_DQ                      (flash_DQ),                                                //                    .export
		.i_avalon_erase_write       (mm_interconnect_0_flash_flash_erase_control_write),       // flash_erase_control.write
		.i_avalon_erase_read        (mm_interconnect_0_flash_flash_erase_control_read),        //                    .read
		.i_avalon_erase_byteenable  (mm_interconnect_0_flash_flash_erase_control_byteenable),  //                    .byteenable
		.i_avalon_erase_writedata   (mm_interconnect_0_flash_flash_erase_control_writedata),   //                    .writedata
		.i_avalon_erase_chip_select (mm_interconnect_0_flash_flash_erase_control_chipselect),  //                    .chipselect
		.o_avalon_erase_readdata    (mm_interconnect_0_flash_flash_erase_control_readdata),    //                    .readdata
		.o_avalon_erase_waitrequest (mm_interconnect_0_flash_flash_erase_control_waitrequest)  //                    .waitrequest
	);

	Computer_System_Green_LEDs green_leds (
		.clk        (system_pll_sys_clk_clk),                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_green_leds_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_green_leds_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_green_leds_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_green_leds_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_green_leds_s1_readdata),   //                    .readdata
		.out_port   (green_leds_export)                           // external_connection.export
	);

	Computer_System_HEX3_HEX0 hex3_hex0 (
		.clk        (system_pll_sys_clk_clk),                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_hex3_hex0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex3_hex0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex3_hex0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex3_hex0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex3_hex0_s1_readdata),   //                    .readdata
		.out_port   (hex3_hex0_export)                           // external_connection.export
	);

	Computer_System_HEX3_HEX0 hex7_hex4 (
		.clk        (system_pll_sys_clk_clk),                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_hex7_hex4_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex7_hex4_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex7_hex4_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex7_hex4_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex7_hex4_s1_readdata),   //                    .readdata
		.out_port   (hex7_hex4_export)                           // external_connection.export
	);

	Computer_System_Interval_Timer interval_timer (
		.clk        (system_pll_sys_clk_clk),                         //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                // reset.reset_n
		.address    (mm_interconnect_0_interval_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_interval_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_interval_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_interval_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_interval_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver9_irq)                        //   irq.irq
	);

	Computer_System_Interval_Timer interval_timer_2 (
		.clk        (system_pll_sys_clk_clk),                           //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                  // reset.reset_n
		.address    (mm_interconnect_0_interval_timer_2_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_interval_timer_2_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_interval_timer_2_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_interval_timer_2_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_interval_timer_2_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver10_irq)                         //   irq.irq
	);

	Computer_System_Interval_Timer interval_timer_2nd_core (
		.clk        (system_pll_sys_clk_clk),                                  //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                         // reset.reset_n
		.address    (mm_interconnect_0_interval_timer_2nd_core_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_interval_timer_2nd_core_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_interval_timer_2nd_core_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_interval_timer_2nd_core_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_interval_timer_2nd_core_s1_write),     //      .write_n
		.irq        (irq_mapper_001_receiver9_irq)                             //   irq.irq
	);

	Computer_System_Interval_Timer interval_timer_2nd_core_2 (
		.clk        (system_pll_sys_clk_clk),                                    //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                           // reset.reset_n
		.address    (mm_interconnect_0_interval_timer_2nd_core_2_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_interval_timer_2nd_core_2_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_interval_timer_2nd_core_2_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_interval_timer_2nd_core_2_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_interval_timer_2nd_core_2_s1_write),     //      .write_n
		.irq        (irq_mapper_001_receiver10_irq)                              //   irq.irq
	);

	Computer_System_IrDA irda (
		.clk        (system_pll_sys_clk_clk),                              //                clk.clk
		.reset      (rst_controller_reset_out_reset),                      //              reset.reset
		.address    (mm_interconnect_0_irda_avalon_irda_slave_address),    //  avalon_irda_slave.address
		.chipselect (mm_interconnect_0_irda_avalon_irda_slave_chipselect), //                   .chipselect
		.byteenable (mm_interconnect_0_irda_avalon_irda_slave_byteenable), //                   .byteenable
		.read       (mm_interconnect_0_irda_avalon_irda_slave_read),       //                   .read
		.write      (mm_interconnect_0_irda_avalon_irda_slave_write),      //                   .write
		.writedata  (mm_interconnect_0_irda_avalon_irda_slave_writedata),  //                   .writedata
		.readdata   (mm_interconnect_0_irda_avalon_irda_slave_readdata),   //                   .readdata
		.irq        (irq_mapper_receiver5_irq),                            //          interrupt.irq
		.IRDA_TXD   (irda_TXD),                                            // external_interface.export
		.IRDA_RXD   (irda_RXD)                                             //                   .export
	);

	Computer_System_JTAG_UART jtag_uart (
		.clk            (system_pll_sys_clk_clk),                                    //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver8_irq)                                   //               irq.irq
	);

	Computer_System_JTAG_UART jtag_uart_2nd_core (
		.clk            (system_pll_sys_clk_clk),                                             //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                                    //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_001_receiver8_irq)                                        //               irq.irq
	);

	Computer_System_JTAG_to_FPGA_Bridge #(
		.USE_PLI     (0),
		.PLI_PORT    (50000),
		.FIFO_DEPTHS (2)
	) jtag_to_fpga_bridge (
		.clk_clk              (system_pll_sys_clk_clk),                   //          clk.clk
		.clk_reset_reset      (system_pll_reset_source_reset),            //    clk_reset.reset
		.master_address       (jtag_to_fpga_bridge_master_address),       //       master.address
		.master_readdata      (jtag_to_fpga_bridge_master_readdata),      //             .readdata
		.master_read          (jtag_to_fpga_bridge_master_read),          //             .read
		.master_write         (jtag_to_fpga_bridge_master_write),         //             .write
		.master_writedata     (jtag_to_fpga_bridge_master_writedata),     //             .writedata
		.master_waitrequest   (jtag_to_fpga_bridge_master_waitrequest),   //             .waitrequest
		.master_readdatavalid (jtag_to_fpga_bridge_master_readdatavalid), //             .readdatavalid
		.master_byteenable    (jtag_to_fpga_bridge_master_byteenable),    //             .byteenable
		.master_reset_reset   ()                                          // master_reset.reset
	);

	Computer_System_Nios2 nios2 (
		.clk                                 (system_pll_sys_clk_clk),                              //                       clk.clk
		.reset_n                             (~rst_controller_001_reset_out_reset),                 //                     reset.reset_n
		.d_address                           (nios2_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_data_master_read),                              //                          .read
		.d_readdata                          (nios2_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_data_master_write),                             //                          .write
		.d_writedata                         (nios2_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (nios2_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (nios2_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_debug_mem_slave_writedata),   //                          .writedata
		.A_ci_multi_done                     (nios2_custom_instruction_master_done),                // custom_instruction_master.done
		.A_ci_multi_result                   (nios2_custom_instruction_master_multi_result),        //                          .multi_result
		.A_ci_multi_a                        (nios2_custom_instruction_master_multi_a),             //                          .multi_a
		.A_ci_multi_b                        (nios2_custom_instruction_master_multi_b),             //                          .multi_b
		.A_ci_multi_c                        (nios2_custom_instruction_master_multi_c),             //                          .multi_c
		.A_ci_multi_clk_en                   (nios2_custom_instruction_master_clk_en),              //                          .clk_en
		.A_ci_multi_clock                    (nios2_custom_instruction_master_clk),                 //                          .clk
		.A_ci_multi_reset                    (nios2_custom_instruction_master_reset),               //                          .reset
		.A_ci_multi_reset_req                (nios2_custom_instruction_master_reset_req),           //                          .reset_req
		.A_ci_multi_dataa                    (nios2_custom_instruction_master_multi_dataa),         //                          .multi_dataa
		.A_ci_multi_datab                    (nios2_custom_instruction_master_multi_datab),         //                          .multi_datab
		.A_ci_multi_n                        (nios2_custom_instruction_master_multi_n),             //                          .multi_n
		.A_ci_multi_readra                   (nios2_custom_instruction_master_multi_readra),        //                          .multi_readra
		.A_ci_multi_readrb                   (nios2_custom_instruction_master_multi_readrb),        //                          .multi_readrb
		.A_ci_multi_start                    (nios2_custom_instruction_master_start),               //                          .start
		.A_ci_multi_writerc                  (nios2_custom_instruction_master_multi_writerc)        //                          .multi_writerc
	);

	Computer_System_Nios2_2nd_Core nios2_2nd_core (
		.clk                                 (system_pll_sys_clk_clk),                                       //                       clk.clk
		.reset_n                             (~rst_controller_002_reset_out_reset),                          //                     reset.reset_n
		.d_address                           (nios2_2nd_core_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_2nd_core_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_2nd_core_data_master_read),                              //                          .read
		.d_readdata                          (nios2_2nd_core_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_2nd_core_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_2nd_core_data_master_write),                             //                          .write
		.d_writedata                         (nios2_2nd_core_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_2nd_core_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_2nd_core_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_2nd_core_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_2nd_core_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_2nd_core_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (nios2_2nd_core_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (nios2_2nd_core_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_2nd_core_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_2nd_core_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_2nd_core_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_2nd_core_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_2nd_core_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_2nd_core_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_2nd_core_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_2nd_core_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_2nd_core_debug_mem_slave_writedata),   //                          .writedata
		.A_ci_multi_done                     (nios2_2nd_core_custom_instruction_master_done),                // custom_instruction_master.done
		.A_ci_multi_result                   (nios2_2nd_core_custom_instruction_master_multi_result),        //                          .multi_result
		.A_ci_multi_a                        (nios2_2nd_core_custom_instruction_master_multi_a),             //                          .multi_a
		.A_ci_multi_b                        (nios2_2nd_core_custom_instruction_master_multi_b),             //                          .multi_b
		.A_ci_multi_c                        (nios2_2nd_core_custom_instruction_master_multi_c),             //                          .multi_c
		.A_ci_multi_clk_en                   (nios2_2nd_core_custom_instruction_master_clk_en),              //                          .clk_en
		.A_ci_multi_clock                    (nios2_2nd_core_custom_instruction_master_clk),                 //                          .clk
		.A_ci_multi_reset                    (nios2_2nd_core_custom_instruction_master_reset),               //                          .reset
		.A_ci_multi_reset_req                (nios2_2nd_core_custom_instruction_master_reset_req),           //                          .reset_req
		.A_ci_multi_dataa                    (nios2_2nd_core_custom_instruction_master_multi_dataa),         //                          .multi_dataa
		.A_ci_multi_datab                    (nios2_2nd_core_custom_instruction_master_multi_datab),         //                          .multi_datab
		.A_ci_multi_n                        (nios2_2nd_core_custom_instruction_master_multi_n),             //                          .multi_n
		.A_ci_multi_readra                   (nios2_2nd_core_custom_instruction_master_multi_readra),        //                          .multi_readra
		.A_ci_multi_readrb                   (nios2_2nd_core_custom_instruction_master_multi_readrb),        //                          .multi_readrb
		.A_ci_multi_start                    (nios2_2nd_core_custom_instruction_master_start),               //                          .start
		.A_ci_multi_writerc                  (nios2_2nd_core_custom_instruction_master_multi_writerc)        //                          .multi_writerc
	);

	fpoint_wrapper #(
		.useDivider (1)
	) nios2_2nd_core_floating_point (
		.clk    (nios2_2nd_core_custom_instruction_master_multi_slave_translator0_ci_master_clk),    // s1.clk
		.clk_en (nios2_2nd_core_custom_instruction_master_multi_slave_translator0_ci_master_clk_en), //   .clk_en
		.dataa  (nios2_2nd_core_custom_instruction_master_multi_slave_translator0_ci_master_dataa),  //   .dataa
		.datab  (nios2_2nd_core_custom_instruction_master_multi_slave_translator0_ci_master_datab),  //   .datab
		.n      (nios2_2nd_core_custom_instruction_master_multi_slave_translator0_ci_master_n),      //   .n
		.reset  (nios2_2nd_core_custom_instruction_master_multi_slave_translator0_ci_master_reset),  //   .reset
		.start  (nios2_2nd_core_custom_instruction_master_multi_slave_translator0_ci_master_start),  //   .start
		.done   (nios2_2nd_core_custom_instruction_master_multi_slave_translator0_ci_master_done),   //   .done
		.result (nios2_2nd_core_custom_instruction_master_multi_slave_translator0_ci_master_result)  //   .result
	);

	fpoint_wrapper #(
		.useDivider (1)
	) nios2_floating_point (
		.clk    (nios2_custom_instruction_master_multi_slave_translator0_ci_master_clk),    // s1.clk
		.clk_en (nios2_custom_instruction_master_multi_slave_translator0_ci_master_clk_en), //   .clk_en
		.dataa  (nios2_custom_instruction_master_multi_slave_translator0_ci_master_dataa),  //   .dataa
		.datab  (nios2_custom_instruction_master_multi_slave_translator0_ci_master_datab),  //   .datab
		.n      (nios2_custom_instruction_master_multi_slave_translator0_ci_master_n),      //   .n
		.reset  (nios2_custom_instruction_master_multi_slave_translator0_ci_master_reset),  //   .reset
		.start  (nios2_custom_instruction_master_multi_slave_translator0_ci_master_start),  //   .start
		.done   (nios2_custom_instruction_master_multi_slave_translator0_ci_master_done),   //   .done
		.result (nios2_custom_instruction_master_multi_slave_translator0_ci_master_result)  //   .result
	);

	Computer_System_PS2_Port ps2_port (
		.clk         (system_pll_sys_clk_clk),                                  //                clk.clk
		.reset       (rst_controller_reset_out_reset),                          //              reset.reset
		.address     (mm_interconnect_0_ps2_port_avalon_ps2_slave_address),     //   avalon_ps2_slave.address
		.chipselect  (mm_interconnect_0_ps2_port_avalon_ps2_slave_chipselect),  //                   .chipselect
		.byteenable  (mm_interconnect_0_ps2_port_avalon_ps2_slave_byteenable),  //                   .byteenable
		.read        (mm_interconnect_0_ps2_port_avalon_ps2_slave_read),        //                   .read
		.write       (mm_interconnect_0_ps2_port_avalon_ps2_slave_write),       //                   .write
		.writedata   (mm_interconnect_0_ps2_port_avalon_ps2_slave_writedata),   //                   .writedata
		.readdata    (mm_interconnect_0_ps2_port_avalon_ps2_slave_readdata),    //                   .readdata
		.waitrequest (mm_interconnect_0_ps2_port_avalon_ps2_slave_waitrequest), //                   .waitrequest
		.irq         (irq_mapper_receiver1_irq),                                //          interrupt.irq
		.PS2_CLK     (ps2_port_CLK),                                            // external_interface.export
		.PS2_DAT     (ps2_port_DAT)                                             //                   .export
	);

	Computer_System_PS2_Port ps2_port_dual (
		.clk         (system_pll_sys_clk_clk),                                       //                clk.clk
		.reset       (rst_controller_reset_out_reset),                               //              reset.reset
		.address     (mm_interconnect_0_ps2_port_dual_avalon_ps2_slave_address),     //   avalon_ps2_slave.address
		.chipselect  (mm_interconnect_0_ps2_port_dual_avalon_ps2_slave_chipselect),  //                   .chipselect
		.byteenable  (mm_interconnect_0_ps2_port_dual_avalon_ps2_slave_byteenable),  //                   .byteenable
		.read        (mm_interconnect_0_ps2_port_dual_avalon_ps2_slave_read),        //                   .read
		.write       (mm_interconnect_0_ps2_port_dual_avalon_ps2_slave_write),       //                   .write
		.writedata   (mm_interconnect_0_ps2_port_dual_avalon_ps2_slave_writedata),   //                   .writedata
		.readdata    (mm_interconnect_0_ps2_port_dual_avalon_ps2_slave_readdata),    //                   .readdata
		.waitrequest (mm_interconnect_0_ps2_port_dual_avalon_ps2_slave_waitrequest), //                   .waitrequest
		.irq         (irq_mapper_receiver2_irq),                                     //          interrupt.irq
		.PS2_CLK     (ps2_port_dual_CLK),                                            // external_interface.export
		.PS2_DAT     (ps2_port_dual_DAT)                                             //                   .export
	);

	Computer_System_Pushbuttons pushbuttons (
		.clk        (system_pll_sys_clk_clk),                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_pushbuttons_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pushbuttons_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pushbuttons_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pushbuttons_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pushbuttons_s1_readdata),   //                    .readdata
		.in_port    (pushbuttons_export),                          // external_connection.export
		.irq        (irq_mapper_receiver6_irq)                     //                 irq.irq
	);

	Computer_System_Red_LEDs red_leds (
		.clk        (system_pll_sys_clk_clk),                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_red_leds_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_red_leds_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_red_leds_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_red_leds_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_red_leds_s1_readdata),   //                    .readdata
		.out_port   (red_leds_export)                           // external_connection.export
	);

	Computer_System_SDRAM sdram (
		.clk            (system_pll_sys_clk_clk),                   //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),          // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_addr),                               //  wire.export
		.zs_ba          (sdram_ba),                                 //      .export
		.zs_cas_n       (sdram_cas_n),                              //      .export
		.zs_cke         (sdram_cke),                                //      .export
		.zs_cs_n        (sdram_cs_n),                               //      .export
		.zs_dq          (sdram_dq),                                 //      .export
		.zs_dqm         (sdram_dqm),                                //      .export
		.zs_ras_n       (sdram_ras_n),                              //      .export
		.zs_we_n        (sdram_we_n)                                //      .export
	);

	Altera_UP_SD_Card_Avalon_Interface sd_card (
		.i_avalon_chip_select (mm_interconnect_0_sd_card_avalon_sdcard_slave_chipselect),  // avalon_sdcard_slave.chipselect
		.i_avalon_address     (mm_interconnect_0_sd_card_avalon_sdcard_slave_address),     //                    .address
		.i_avalon_read        (mm_interconnect_0_sd_card_avalon_sdcard_slave_read),        //                    .read
		.i_avalon_write       (mm_interconnect_0_sd_card_avalon_sdcard_slave_write),       //                    .write
		.i_avalon_byteenable  (mm_interconnect_0_sd_card_avalon_sdcard_slave_byteenable),  //                    .byteenable
		.i_avalon_writedata   (mm_interconnect_0_sd_card_avalon_sdcard_slave_writedata),   //                    .writedata
		.o_avalon_readdata    (mm_interconnect_0_sd_card_avalon_sdcard_slave_readdata),    //                    .readdata
		.o_avalon_waitrequest (mm_interconnect_0_sd_card_avalon_sdcard_slave_waitrequest), //                    .waitrequest
		.i_clock              (system_pll_sys_clk_clk),                                    //                 clk.clk
		.i_reset_n            (~rst_controller_reset_out_reset),                           //               reset.reset_n
		.b_SD_cmd             (sd_card_b_SD_cmd),                                          //         conduit_end.export
		.b_SD_dat             (sd_card_b_SD_dat),                                          //                    .export
		.b_SD_dat3            (sd_card_b_SD_dat3),                                         //                    .export
		.o_SD_clock           (sd_card_o_SD_clock)                                         //                    .export
	);

	Computer_System_SRAM sram (
		.clk           (system_pll_sys_clk_clk),                                 //                clk.clk
		.reset         (rst_controller_reset_out_reset),                         //              reset.reset
		.SRAM_DQ       (sram_DQ),                                                // external_interface.export
		.SRAM_ADDR     (sram_ADDR),                                              //                   .export
		.SRAM_LB_N     (sram_LB_N),                                              //                   .export
		.SRAM_UB_N     (sram_UB_N),                                              //                   .export
		.SRAM_CE_N     (sram_CE_N),                                              //                   .export
		.SRAM_OE_N     (sram_OE_N),                                              //                   .export
		.SRAM_WE_N     (sram_WE_N),                                              //                   .export
		.address       (mm_interconnect_0_sram_avalon_sram_slave_address),       //  avalon_sram_slave.address
		.byteenable    (mm_interconnect_0_sram_avalon_sram_slave_byteenable),    //                   .byteenable
		.read          (mm_interconnect_0_sram_avalon_sram_slave_read),          //                   .read
		.write         (mm_interconnect_0_sram_avalon_sram_slave_write),         //                   .write
		.writedata     (mm_interconnect_0_sram_avalon_sram_slave_writedata),     //                   .writedata
		.readdata      (mm_interconnect_0_sram_avalon_sram_slave_readdata),      //                   .readdata
		.readdatavalid (mm_interconnect_0_sram_avalon_sram_slave_readdatavalid)  //                   .readdatavalid
	);

	Computer_System_Serial_Port serial_port (
		.clk        (system_pll_sys_clk_clk),                                      //                clk.clk
		.reset      (rst_controller_reset_out_reset),                              //              reset.reset
		.address    (mm_interconnect_0_serial_port_avalon_rs232_slave_address),    // avalon_rs232_slave.address
		.chipselect (mm_interconnect_0_serial_port_avalon_rs232_slave_chipselect), //                   .chipselect
		.byteenable (mm_interconnect_0_serial_port_avalon_rs232_slave_byteenable), //                   .byteenable
		.read       (mm_interconnect_0_serial_port_avalon_rs232_slave_read),       //                   .read
		.write      (mm_interconnect_0_serial_port_avalon_rs232_slave_write),      //                   .write
		.writedata  (mm_interconnect_0_serial_port_avalon_rs232_slave_writedata),  //                   .writedata
		.readdata   (mm_interconnect_0_serial_port_avalon_rs232_slave_readdata),   //                   .readdata
		.irq        (irq_mapper_receiver4_irq),                                    //          interrupt.irq
		.UART_RXD   (serial_port_RXD),                                             // external_interface.export
		.UART_TXD   (serial_port_TXD)                                              //                   .export
	);

	Computer_System_Slider_Switches slider_switches (
		.clk      (system_pll_sys_clk_clk),                        //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address  (mm_interconnect_0_slider_switches_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_slider_switches_s1_readdata), //                    .readdata
		.in_port  (slider_switches_export)                         // external_connection.export
	);

	Computer_System_SysID sysid (
		.clock    (system_pll_sys_clk_clk),                         //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_control_slave_address)   //              .address
	);

	Computer_System_System_PLL system_pll (
		.ref_clk_clk        (system_pll_ref_clk_clk),        //      ref_clk.clk
		.ref_reset_reset    (system_pll_ref_reset_reset),    //    ref_reset.reset
		.sys_clk_clk        (system_pll_sys_clk_clk),        //      sys_clk.clk
		.sdram_clk_clk      (sdram_clk_clk),                 //    sdram_clk.clk
		.reset_source_reset (system_pll_reset_source_reset)  // reset_source.reset
	);

	Computer_System_USB usb (
		.clk        (system_pll_sys_clk_clk),                            //                clk.clk
		.reset      (rst_controller_reset_out_reset),                    //              reset.reset
		.address    (mm_interconnect_0_usb_avalon_usb_slave_address),    //   avalon_usb_slave.address
		.chipselect (mm_interconnect_0_usb_avalon_usb_slave_chipselect), //                   .chipselect
		.read       (mm_interconnect_0_usb_avalon_usb_slave_read),       //                   .read
		.write      (mm_interconnect_0_usb_avalon_usb_slave_write),      //                   .write
		.writedata  (mm_interconnect_0_usb_avalon_usb_slave_writedata),  //                   .writedata
		.readdata   (mm_interconnect_0_usb_avalon_usb_slave_readdata),   //                   .readdata
		.irq        (irq_mapper_receiver3_irq),                          //          interrupt.irq
		.OTG_INT1   (usb_INT1),                                          // external_interface.export
		.OTG_DATA   (usb_DATA),                                          //                   .export
		.OTG_RST_N  (usb_RST_N),                                         //                   .export
		.OTG_ADDR   (usb_ADDR),                                          //                   .export
		.OTG_CS_N   (usb_CS_N),                                          //                   .export
		.OTG_RD_N   (usb_RD_N),                                          //                   .export
		.OTG_WR_N   (usb_WR_N),                                          //                   .export
		.OTG_INT0   (usb_INT0)                                           //                   .export
	);

	Computer_System_VGA_Subsystem vga_subsystem (
		.char_buffer_control_slave_address    (mm_interconnect_0_vga_subsystem_char_buffer_control_slave_address),    // char_buffer_control_slave.address
		.char_buffer_control_slave_byteenable (mm_interconnect_0_vga_subsystem_char_buffer_control_slave_byteenable), //                          .byteenable
		.char_buffer_control_slave_read       (mm_interconnect_0_vga_subsystem_char_buffer_control_slave_read),       //                          .read
		.char_buffer_control_slave_write      (mm_interconnect_0_vga_subsystem_char_buffer_control_slave_write),      //                          .write
		.char_buffer_control_slave_writedata  (mm_interconnect_0_vga_subsystem_char_buffer_control_slave_writedata),  //                          .writedata
		.char_buffer_control_slave_readdata   (mm_interconnect_0_vga_subsystem_char_buffer_control_slave_readdata),   //                          .readdata
		.char_buffer_slave_address            (mm_interconnect_0_vga_subsystem_char_buffer_slave_address),            //         char_buffer_slave.address
		.char_buffer_slave_clken              (mm_interconnect_0_vga_subsystem_char_buffer_slave_clken),              //                          .clken
		.char_buffer_slave_chipselect         (mm_interconnect_0_vga_subsystem_char_buffer_slave_chipselect),         //                          .chipselect
		.char_buffer_slave_write              (mm_interconnect_0_vga_subsystem_char_buffer_slave_write),              //                          .write
		.char_buffer_slave_readdata           (mm_interconnect_0_vga_subsystem_char_buffer_slave_readdata),           //                          .readdata
		.char_buffer_slave_writedata          (mm_interconnect_0_vga_subsystem_char_buffer_slave_writedata),          //                          .writedata
		.char_buffer_slave_byteenable         (mm_interconnect_0_vga_subsystem_char_buffer_slave_byteenable),         //                          .byteenable
		.pixel_dma_control_slave_address      (mm_interconnect_0_vga_subsystem_pixel_dma_control_slave_address),      //   pixel_dma_control_slave.address
		.pixel_dma_control_slave_byteenable   (mm_interconnect_0_vga_subsystem_pixel_dma_control_slave_byteenable),   //                          .byteenable
		.pixel_dma_control_slave_read         (mm_interconnect_0_vga_subsystem_pixel_dma_control_slave_read),         //                          .read
		.pixel_dma_control_slave_write        (mm_interconnect_0_vga_subsystem_pixel_dma_control_slave_write),        //                          .write
		.pixel_dma_control_slave_writedata    (mm_interconnect_0_vga_subsystem_pixel_dma_control_slave_writedata),    //                          .writedata
		.pixel_dma_control_slave_readdata     (mm_interconnect_0_vga_subsystem_pixel_dma_control_slave_readdata),     //                          .readdata
		.pixel_dma_master_address             (vga_subsystem_pixel_dma_master_address),                               //          pixel_dma_master.address
		.pixel_dma_master_waitrequest         (vga_subsystem_pixel_dma_master_waitrequest),                           //                          .waitrequest
		.pixel_dma_master_lock                (vga_subsystem_pixel_dma_master_lock),                                  //                          .lock
		.pixel_dma_master_read                (vga_subsystem_pixel_dma_master_read),                                  //                          .read
		.pixel_dma_master_readdata            (vga_subsystem_pixel_dma_master_readdata),                              //                          .readdata
		.pixel_dma_master_readdatavalid       (vga_subsystem_pixel_dma_master_readdatavalid),                         //                          .readdatavalid
		.rgb_slave_read                       (mm_interconnect_0_vga_subsystem_rgb_slave_read),                       //                 rgb_slave.read
		.rgb_slave_readdata                   (mm_interconnect_0_vga_subsystem_rgb_slave_readdata),                   //                          .readdata
		.sys_clk_clk                          (system_pll_sys_clk_clk),                                               //                   sys_clk.clk
		.sys_reset_reset_n                    (~system_pll_reset_source_reset),                                       //                 sys_reset.reset_n
		.vga_CLK                              (vga_CLK),                                                              //                       vga.CLK
		.vga_HS                               (vga_HS),                                                               //                          .HS
		.vga_VS                               (vga_VS),                                                               //                          .VS
		.vga_BLANK                            (vga_BLANK),                                                            //                          .BLANK
		.vga_SYNC                             (vga_SYNC),                                                             //                          .SYNC
		.vga_R                                (vga_R),                                                                //                          .R
		.vga_G                                (vga_G),                                                                //                          .G
		.vga_B                                (vga_B),                                                                //                          .B
		.vga_clk_clk                          (video_pll_vga_clk_clk),                                                //                   vga_clk.clk
		.vga_reset_reset_n                    (~video_pll_reset_source_reset)                                         //                 vga_reset.reset_n
	);

	Computer_System_Video_In_Subsystem video_in_subsystem (
		.sys_clk_clk                                      (system_pll_sys_clk_clk),                                                                //                               sys_clk.clk
		.sys_reset_reset_n                                (~system_pll_reset_source_reset),                                                        //                             sys_reset.reset_n
		.video_in_TD_CLK27                                (video_in_TD_CLK27),                                                                     //                              video_in.TD_CLK27
		.video_in_TD_DATA                                 (video_in_TD_DATA),                                                                      //                                      .TD_DATA
		.video_in_TD_HS                                   (video_in_TD_HS),                                                                        //                                      .TD_HS
		.video_in_TD_VS                                   (video_in_TD_VS),                                                                        //                                      .TD_VS
		.video_in_clk27_reset                             (video_in_clk27_reset),                                                                  //                                      .clk27_reset
		.video_in_TD_RESET                                (video_in_TD_RESET),                                                                     //                                      .TD_RESET
		.video_in_overflow_flag                           (video_in_overflow_flag),                                                                //                                      .overflow_flag
		.video_in_dma_control_slave_address               (mm_interconnect_0_video_in_subsystem_video_in_dma_control_slave_address),               //            video_in_dma_control_slave.address
		.video_in_dma_control_slave_byteenable            (mm_interconnect_0_video_in_subsystem_video_in_dma_control_slave_byteenable),            //                                      .byteenable
		.video_in_dma_control_slave_read                  (mm_interconnect_0_video_in_subsystem_video_in_dma_control_slave_read),                  //                                      .read
		.video_in_dma_control_slave_write                 (mm_interconnect_0_video_in_subsystem_video_in_dma_control_slave_write),                 //                                      .write
		.video_in_dma_control_slave_writedata             (mm_interconnect_0_video_in_subsystem_video_in_dma_control_slave_writedata),             //                                      .writedata
		.video_in_dma_control_slave_readdata              (mm_interconnect_0_video_in_subsystem_video_in_dma_control_slave_readdata),              //                                      .readdata
		.video_in_dma_master_address                      (video_in_subsystem_video_in_dma_master_address),                                        //                   video_in_dma_master.address
		.video_in_dma_master_waitrequest                  (video_in_subsystem_video_in_dma_master_waitrequest),                                    //                                      .waitrequest
		.video_in_dma_master_write                        (video_in_subsystem_video_in_dma_master_write),                                          //                                      .write
		.video_in_dma_master_writedata                    (video_in_subsystem_video_in_dma_master_writedata),                                      //                                      .writedata
		.video_in_edge_detection_control_slave_address    (mm_interconnect_0_video_in_subsystem_video_in_edge_detection_control_slave_address),    // video_in_edge_detection_control_slave.address
		.video_in_edge_detection_control_slave_write_n    (~mm_interconnect_0_video_in_subsystem_video_in_edge_detection_control_slave_write),     //                                      .write_n
		.video_in_edge_detection_control_slave_writedata  (mm_interconnect_0_video_in_subsystem_video_in_edge_detection_control_slave_writedata),  //                                      .writedata
		.video_in_edge_detection_control_slave_chipselect (mm_interconnect_0_video_in_subsystem_video_in_edge_detection_control_slave_chipselect), //                                      .chipselect
		.video_in_edge_detection_control_slave_readdata   (mm_interconnect_0_video_in_subsystem_video_in_edge_detection_control_slave_readdata)    //                                      .readdata
	);

	Computer_System_Video_PLL video_pll (
		.ref_clk_clk        (video_pll_ref_clk_clk),        //      ref_clk.clk
		.ref_reset_reset    (video_pll_ref_reset_reset),    //    ref_reset.reset
		.vga_clk_clk        (video_pll_vga_clk_clk),        //      vga_clk.clk
		.reset_source_reset (video_pll_reset_source_reset)  // reset_source.reset
	);

	gcd_ci hw_convolution_inst_0 (
		.clk_en (nios2_custom_instruction_master_multi_slave_translator1_ci_master_clk_en), // nios_custom_instruction_slave.clk_en
		.dataa  (nios2_custom_instruction_master_multi_slave_translator1_ci_master_dataa),  //                              .dataa
		.datab  (nios2_custom_instruction_master_multi_slave_translator1_ci_master_datab),  //                              .datab
		.result (nios2_custom_instruction_master_multi_slave_translator1_ci_master_result), //                              .result
		.start  (nios2_custom_instruction_master_multi_slave_translator1_ci_master_start),  //                              .start
		.done   (nios2_custom_instruction_master_multi_slave_translator1_ci_master_done),   //                              .done
		.clk    (nios2_custom_instruction_master_multi_slave_translator1_ci_master_clk),    //                              .clk
		.reset  (nios2_custom_instruction_master_multi_slave_translator1_ci_master_reset)   //                              .reset
	);

	altera_customins_master_translator #(
		.SHARED_COMB_AND_MULTI (0)
	) nios2_custom_instruction_master_translator (
		.ci_slave_result           (),                                                                     //        ci_slave.result
		.ci_slave_multi_clk        (nios2_custom_instruction_master_clk),                                  //                .clk
		.ci_slave_multi_reset      (nios2_custom_instruction_master_reset),                                //                .reset
		.ci_slave_multi_clken      (nios2_custom_instruction_master_clk_en),                               //                .clk_en
		.ci_slave_multi_reset_req  (nios2_custom_instruction_master_reset_req),                            //                .reset_req
		.ci_slave_multi_start      (nios2_custom_instruction_master_start),                                //                .start
		.ci_slave_multi_done       (nios2_custom_instruction_master_done),                                 //                .done
		.ci_slave_multi_dataa      (nios2_custom_instruction_master_multi_dataa),                          //                .multi_dataa
		.ci_slave_multi_datab      (nios2_custom_instruction_master_multi_datab),                          //                .multi_datab
		.ci_slave_multi_result     (nios2_custom_instruction_master_multi_result),                         //                .multi_result
		.ci_slave_multi_n          (nios2_custom_instruction_master_multi_n),                              //                .multi_n
		.ci_slave_multi_readra     (nios2_custom_instruction_master_multi_readra),                         //                .multi_readra
		.ci_slave_multi_readrb     (nios2_custom_instruction_master_multi_readrb),                         //                .multi_readrb
		.ci_slave_multi_writerc    (nios2_custom_instruction_master_multi_writerc),                        //                .multi_writerc
		.ci_slave_multi_a          (nios2_custom_instruction_master_multi_a),                              //                .multi_a
		.ci_slave_multi_b          (nios2_custom_instruction_master_multi_b),                              //                .multi_b
		.ci_slave_multi_c          (nios2_custom_instruction_master_multi_c),                              //                .multi_c
		.comb_ci_master_result     (),                                                                     //  comb_ci_master.result
		.multi_ci_master_clk       (nios2_custom_instruction_master_translator_multi_ci_master_clk),       // multi_ci_master.clk
		.multi_ci_master_reset     (nios2_custom_instruction_master_translator_multi_ci_master_reset),     //                .reset
		.multi_ci_master_clken     (nios2_custom_instruction_master_translator_multi_ci_master_clk_en),    //                .clk_en
		.multi_ci_master_reset_req (nios2_custom_instruction_master_translator_multi_ci_master_reset_req), //                .reset_req
		.multi_ci_master_start     (nios2_custom_instruction_master_translator_multi_ci_master_start),     //                .start
		.multi_ci_master_done      (nios2_custom_instruction_master_translator_multi_ci_master_done),      //                .done
		.multi_ci_master_dataa     (nios2_custom_instruction_master_translator_multi_ci_master_dataa),     //                .dataa
		.multi_ci_master_datab     (nios2_custom_instruction_master_translator_multi_ci_master_datab),     //                .datab
		.multi_ci_master_result    (nios2_custom_instruction_master_translator_multi_ci_master_result),    //                .result
		.multi_ci_master_n         (nios2_custom_instruction_master_translator_multi_ci_master_n),         //                .n
		.multi_ci_master_readra    (nios2_custom_instruction_master_translator_multi_ci_master_readra),    //                .readra
		.multi_ci_master_readrb    (nios2_custom_instruction_master_translator_multi_ci_master_readrb),    //                .readrb
		.multi_ci_master_writerc   (nios2_custom_instruction_master_translator_multi_ci_master_writerc),   //                .writerc
		.multi_ci_master_a         (nios2_custom_instruction_master_translator_multi_ci_master_a),         //                .a
		.multi_ci_master_b         (nios2_custom_instruction_master_translator_multi_ci_master_b),         //                .b
		.multi_ci_master_c         (nios2_custom_instruction_master_translator_multi_ci_master_c),         //                .c
		.ci_slave_dataa            (32'b00000000000000000000000000000000),                                 //     (terminated)
		.ci_slave_datab            (32'b00000000000000000000000000000000),                                 //     (terminated)
		.ci_slave_n                (8'b00000000),                                                          //     (terminated)
		.ci_slave_readra           (1'b0),                                                                 //     (terminated)
		.ci_slave_readrb           (1'b0),                                                                 //     (terminated)
		.ci_slave_writerc          (1'b0),                                                                 //     (terminated)
		.ci_slave_a                (5'b00000),                                                             //     (terminated)
		.ci_slave_b                (5'b00000),                                                             //     (terminated)
		.ci_slave_c                (5'b00000),                                                             //     (terminated)
		.ci_slave_ipending         (32'b00000000000000000000000000000000),                                 //     (terminated)
		.ci_slave_estatus          (1'b0),                                                                 //     (terminated)
		.comb_ci_master_dataa      (),                                                                     //     (terminated)
		.comb_ci_master_datab      (),                                                                     //     (terminated)
		.comb_ci_master_n          (),                                                                     //     (terminated)
		.comb_ci_master_readra     (),                                                                     //     (terminated)
		.comb_ci_master_readrb     (),                                                                     //     (terminated)
		.comb_ci_master_writerc    (),                                                                     //     (terminated)
		.comb_ci_master_a          (),                                                                     //     (terminated)
		.comb_ci_master_b          (),                                                                     //     (terminated)
		.comb_ci_master_c          (),                                                                     //     (terminated)
		.comb_ci_master_ipending   (),                                                                     //     (terminated)
		.comb_ci_master_estatus    ()                                                                      //     (terminated)
	);

	Computer_System_Nios2_custom_instruction_master_multi_xconnect nios2_custom_instruction_master_multi_xconnect (
		.ci_slave_dataa       (nios2_custom_instruction_master_translator_multi_ci_master_dataa),     //   ci_slave.dataa
		.ci_slave_datab       (nios2_custom_instruction_master_translator_multi_ci_master_datab),     //           .datab
		.ci_slave_result      (nios2_custom_instruction_master_translator_multi_ci_master_result),    //           .result
		.ci_slave_n           (nios2_custom_instruction_master_translator_multi_ci_master_n),         //           .n
		.ci_slave_readra      (nios2_custom_instruction_master_translator_multi_ci_master_readra),    //           .readra
		.ci_slave_readrb      (nios2_custom_instruction_master_translator_multi_ci_master_readrb),    //           .readrb
		.ci_slave_writerc     (nios2_custom_instruction_master_translator_multi_ci_master_writerc),   //           .writerc
		.ci_slave_a           (nios2_custom_instruction_master_translator_multi_ci_master_a),         //           .a
		.ci_slave_b           (nios2_custom_instruction_master_translator_multi_ci_master_b),         //           .b
		.ci_slave_c           (nios2_custom_instruction_master_translator_multi_ci_master_c),         //           .c
		.ci_slave_ipending    (),                                                                     //           .ipending
		.ci_slave_estatus     (),                                                                     //           .estatus
		.ci_slave_clk         (nios2_custom_instruction_master_translator_multi_ci_master_clk),       //           .clk
		.ci_slave_reset       (nios2_custom_instruction_master_translator_multi_ci_master_reset),     //           .reset
		.ci_slave_clken       (nios2_custom_instruction_master_translator_multi_ci_master_clk_en),    //           .clk_en
		.ci_slave_reset_req   (nios2_custom_instruction_master_translator_multi_ci_master_reset_req), //           .reset_req
		.ci_slave_start       (nios2_custom_instruction_master_translator_multi_ci_master_start),     //           .start
		.ci_slave_done        (nios2_custom_instruction_master_translator_multi_ci_master_done),      //           .done
		.ci_master0_dataa     (nios2_custom_instruction_master_multi_xconnect_ci_master0_dataa),      // ci_master0.dataa
		.ci_master0_datab     (nios2_custom_instruction_master_multi_xconnect_ci_master0_datab),      //           .datab
		.ci_master0_result    (nios2_custom_instruction_master_multi_xconnect_ci_master0_result),     //           .result
		.ci_master0_n         (nios2_custom_instruction_master_multi_xconnect_ci_master0_n),          //           .n
		.ci_master0_readra    (nios2_custom_instruction_master_multi_xconnect_ci_master0_readra),     //           .readra
		.ci_master0_readrb    (nios2_custom_instruction_master_multi_xconnect_ci_master0_readrb),     //           .readrb
		.ci_master0_writerc   (nios2_custom_instruction_master_multi_xconnect_ci_master0_writerc),    //           .writerc
		.ci_master0_a         (nios2_custom_instruction_master_multi_xconnect_ci_master0_a),          //           .a
		.ci_master0_b         (nios2_custom_instruction_master_multi_xconnect_ci_master0_b),          //           .b
		.ci_master0_c         (nios2_custom_instruction_master_multi_xconnect_ci_master0_c),          //           .c
		.ci_master0_ipending  (nios2_custom_instruction_master_multi_xconnect_ci_master0_ipending),   //           .ipending
		.ci_master0_estatus   (nios2_custom_instruction_master_multi_xconnect_ci_master0_estatus),    //           .estatus
		.ci_master0_clk       (nios2_custom_instruction_master_multi_xconnect_ci_master0_clk),        //           .clk
		.ci_master0_reset     (nios2_custom_instruction_master_multi_xconnect_ci_master0_reset),      //           .reset
		.ci_master0_clken     (nios2_custom_instruction_master_multi_xconnect_ci_master0_clk_en),     //           .clk_en
		.ci_master0_reset_req (nios2_custom_instruction_master_multi_xconnect_ci_master0_reset_req),  //           .reset_req
		.ci_master0_start     (nios2_custom_instruction_master_multi_xconnect_ci_master0_start),      //           .start
		.ci_master0_done      (nios2_custom_instruction_master_multi_xconnect_ci_master0_done),       //           .done
		.ci_master1_dataa     (nios2_custom_instruction_master_multi_xconnect_ci_master1_dataa),      // ci_master1.dataa
		.ci_master1_datab     (nios2_custom_instruction_master_multi_xconnect_ci_master1_datab),      //           .datab
		.ci_master1_result    (nios2_custom_instruction_master_multi_xconnect_ci_master1_result),     //           .result
		.ci_master1_n         (nios2_custom_instruction_master_multi_xconnect_ci_master1_n),          //           .n
		.ci_master1_readra    (nios2_custom_instruction_master_multi_xconnect_ci_master1_readra),     //           .readra
		.ci_master1_readrb    (nios2_custom_instruction_master_multi_xconnect_ci_master1_readrb),     //           .readrb
		.ci_master1_writerc   (nios2_custom_instruction_master_multi_xconnect_ci_master1_writerc),    //           .writerc
		.ci_master1_a         (nios2_custom_instruction_master_multi_xconnect_ci_master1_a),          //           .a
		.ci_master1_b         (nios2_custom_instruction_master_multi_xconnect_ci_master1_b),          //           .b
		.ci_master1_c         (nios2_custom_instruction_master_multi_xconnect_ci_master1_c),          //           .c
		.ci_master1_ipending  (nios2_custom_instruction_master_multi_xconnect_ci_master1_ipending),   //           .ipending
		.ci_master1_estatus   (nios2_custom_instruction_master_multi_xconnect_ci_master1_estatus),    //           .estatus
		.ci_master1_clk       (nios2_custom_instruction_master_multi_xconnect_ci_master1_clk),        //           .clk
		.ci_master1_reset     (nios2_custom_instruction_master_multi_xconnect_ci_master1_reset),      //           .reset
		.ci_master1_clken     (nios2_custom_instruction_master_multi_xconnect_ci_master1_clk_en),     //           .clk_en
		.ci_master1_reset_req (nios2_custom_instruction_master_multi_xconnect_ci_master1_reset_req),  //           .reset_req
		.ci_master1_start     (nios2_custom_instruction_master_multi_xconnect_ci_master1_start),      //           .start
		.ci_master1_done      (nios2_custom_instruction_master_multi_xconnect_ci_master1_done)        //           .done
	);

	altera_customins_slave_translator #(
		.N_WIDTH          (2),
		.USE_DONE         (1),
		.NUM_FIXED_CYCLES (1)
	) nios2_custom_instruction_master_multi_slave_translator0 (
		.ci_slave_dataa      (nios2_custom_instruction_master_multi_xconnect_ci_master0_dataa),          //  ci_slave.dataa
		.ci_slave_datab      (nios2_custom_instruction_master_multi_xconnect_ci_master0_datab),          //          .datab
		.ci_slave_result     (nios2_custom_instruction_master_multi_xconnect_ci_master0_result),         //          .result
		.ci_slave_n          (nios2_custom_instruction_master_multi_xconnect_ci_master0_n),              //          .n
		.ci_slave_readra     (nios2_custom_instruction_master_multi_xconnect_ci_master0_readra),         //          .readra
		.ci_slave_readrb     (nios2_custom_instruction_master_multi_xconnect_ci_master0_readrb),         //          .readrb
		.ci_slave_writerc    (nios2_custom_instruction_master_multi_xconnect_ci_master0_writerc),        //          .writerc
		.ci_slave_a          (nios2_custom_instruction_master_multi_xconnect_ci_master0_a),              //          .a
		.ci_slave_b          (nios2_custom_instruction_master_multi_xconnect_ci_master0_b),              //          .b
		.ci_slave_c          (nios2_custom_instruction_master_multi_xconnect_ci_master0_c),              //          .c
		.ci_slave_ipending   (nios2_custom_instruction_master_multi_xconnect_ci_master0_ipending),       //          .ipending
		.ci_slave_estatus    (nios2_custom_instruction_master_multi_xconnect_ci_master0_estatus),        //          .estatus
		.ci_slave_clk        (nios2_custom_instruction_master_multi_xconnect_ci_master0_clk),            //          .clk
		.ci_slave_clken      (nios2_custom_instruction_master_multi_xconnect_ci_master0_clk_en),         //          .clk_en
		.ci_slave_reset_req  (nios2_custom_instruction_master_multi_xconnect_ci_master0_reset_req),      //          .reset_req
		.ci_slave_reset      (nios2_custom_instruction_master_multi_xconnect_ci_master0_reset),          //          .reset
		.ci_slave_start      (nios2_custom_instruction_master_multi_xconnect_ci_master0_start),          //          .start
		.ci_slave_done       (nios2_custom_instruction_master_multi_xconnect_ci_master0_done),           //          .done
		.ci_master_dataa     (nios2_custom_instruction_master_multi_slave_translator0_ci_master_dataa),  // ci_master.dataa
		.ci_master_datab     (nios2_custom_instruction_master_multi_slave_translator0_ci_master_datab),  //          .datab
		.ci_master_result    (nios2_custom_instruction_master_multi_slave_translator0_ci_master_result), //          .result
		.ci_master_n         (nios2_custom_instruction_master_multi_slave_translator0_ci_master_n),      //          .n
		.ci_master_clk       (nios2_custom_instruction_master_multi_slave_translator0_ci_master_clk),    //          .clk
		.ci_master_clken     (nios2_custom_instruction_master_multi_slave_translator0_ci_master_clk_en), //          .clk_en
		.ci_master_reset     (nios2_custom_instruction_master_multi_slave_translator0_ci_master_reset),  //          .reset
		.ci_master_start     (nios2_custom_instruction_master_multi_slave_translator0_ci_master_start),  //          .start
		.ci_master_done      (nios2_custom_instruction_master_multi_slave_translator0_ci_master_done),   //          .done
		.ci_master_readra    (),                                                                         // (terminated)
		.ci_master_readrb    (),                                                                         // (terminated)
		.ci_master_writerc   (),                                                                         // (terminated)
		.ci_master_a         (),                                                                         // (terminated)
		.ci_master_b         (),                                                                         // (terminated)
		.ci_master_c         (),                                                                         // (terminated)
		.ci_master_ipending  (),                                                                         // (terminated)
		.ci_master_estatus   (),                                                                         // (terminated)
		.ci_master_reset_req ()                                                                          // (terminated)
	);

	altera_customins_slave_translator #(
		.N_WIDTH          (8),
		.USE_DONE         (1),
		.NUM_FIXED_CYCLES (0)
	) nios2_custom_instruction_master_multi_slave_translator1 (
		.ci_slave_dataa      (nios2_custom_instruction_master_multi_xconnect_ci_master1_dataa),          //  ci_slave.dataa
		.ci_slave_datab      (nios2_custom_instruction_master_multi_xconnect_ci_master1_datab),          //          .datab
		.ci_slave_result     (nios2_custom_instruction_master_multi_xconnect_ci_master1_result),         //          .result
		.ci_slave_n          (nios2_custom_instruction_master_multi_xconnect_ci_master1_n),              //          .n
		.ci_slave_readra     (nios2_custom_instruction_master_multi_xconnect_ci_master1_readra),         //          .readra
		.ci_slave_readrb     (nios2_custom_instruction_master_multi_xconnect_ci_master1_readrb),         //          .readrb
		.ci_slave_writerc    (nios2_custom_instruction_master_multi_xconnect_ci_master1_writerc),        //          .writerc
		.ci_slave_a          (nios2_custom_instruction_master_multi_xconnect_ci_master1_a),              //          .a
		.ci_slave_b          (nios2_custom_instruction_master_multi_xconnect_ci_master1_b),              //          .b
		.ci_slave_c          (nios2_custom_instruction_master_multi_xconnect_ci_master1_c),              //          .c
		.ci_slave_ipending   (nios2_custom_instruction_master_multi_xconnect_ci_master1_ipending),       //          .ipending
		.ci_slave_estatus    (nios2_custom_instruction_master_multi_xconnect_ci_master1_estatus),        //          .estatus
		.ci_slave_clk        (nios2_custom_instruction_master_multi_xconnect_ci_master1_clk),            //          .clk
		.ci_slave_clken      (nios2_custom_instruction_master_multi_xconnect_ci_master1_clk_en),         //          .clk_en
		.ci_slave_reset_req  (nios2_custom_instruction_master_multi_xconnect_ci_master1_reset_req),      //          .reset_req
		.ci_slave_reset      (nios2_custom_instruction_master_multi_xconnect_ci_master1_reset),          //          .reset
		.ci_slave_start      (nios2_custom_instruction_master_multi_xconnect_ci_master1_start),          //          .start
		.ci_slave_done       (nios2_custom_instruction_master_multi_xconnect_ci_master1_done),           //          .done
		.ci_master_dataa     (nios2_custom_instruction_master_multi_slave_translator1_ci_master_dataa),  // ci_master.dataa
		.ci_master_datab     (nios2_custom_instruction_master_multi_slave_translator1_ci_master_datab),  //          .datab
		.ci_master_result    (nios2_custom_instruction_master_multi_slave_translator1_ci_master_result), //          .result
		.ci_master_clk       (nios2_custom_instruction_master_multi_slave_translator1_ci_master_clk),    //          .clk
		.ci_master_clken     (nios2_custom_instruction_master_multi_slave_translator1_ci_master_clk_en), //          .clk_en
		.ci_master_reset     (nios2_custom_instruction_master_multi_slave_translator1_ci_master_reset),  //          .reset
		.ci_master_start     (nios2_custom_instruction_master_multi_slave_translator1_ci_master_start),  //          .start
		.ci_master_done      (nios2_custom_instruction_master_multi_slave_translator1_ci_master_done),   //          .done
		.ci_master_n         (),                                                                         // (terminated)
		.ci_master_readra    (),                                                                         // (terminated)
		.ci_master_readrb    (),                                                                         // (terminated)
		.ci_master_writerc   (),                                                                         // (terminated)
		.ci_master_a         (),                                                                         // (terminated)
		.ci_master_b         (),                                                                         // (terminated)
		.ci_master_c         (),                                                                         // (terminated)
		.ci_master_ipending  (),                                                                         // (terminated)
		.ci_master_estatus   (),                                                                         // (terminated)
		.ci_master_reset_req ()                                                                          // (terminated)
	);

	altera_customins_master_translator #(
		.SHARED_COMB_AND_MULTI (0)
	) nios2_2nd_core_custom_instruction_master_translator (
		.ci_slave_result           (),                                                                              //        ci_slave.result
		.ci_slave_multi_clk        (nios2_2nd_core_custom_instruction_master_clk),                                  //                .clk
		.ci_slave_multi_reset      (nios2_2nd_core_custom_instruction_master_reset),                                //                .reset
		.ci_slave_multi_clken      (nios2_2nd_core_custom_instruction_master_clk_en),                               //                .clk_en
		.ci_slave_multi_reset_req  (nios2_2nd_core_custom_instruction_master_reset_req),                            //                .reset_req
		.ci_slave_multi_start      (nios2_2nd_core_custom_instruction_master_start),                                //                .start
		.ci_slave_multi_done       (nios2_2nd_core_custom_instruction_master_done),                                 //                .done
		.ci_slave_multi_dataa      (nios2_2nd_core_custom_instruction_master_multi_dataa),                          //                .multi_dataa
		.ci_slave_multi_datab      (nios2_2nd_core_custom_instruction_master_multi_datab),                          //                .multi_datab
		.ci_slave_multi_result     (nios2_2nd_core_custom_instruction_master_multi_result),                         //                .multi_result
		.ci_slave_multi_n          (nios2_2nd_core_custom_instruction_master_multi_n),                              //                .multi_n
		.ci_slave_multi_readra     (nios2_2nd_core_custom_instruction_master_multi_readra),                         //                .multi_readra
		.ci_slave_multi_readrb     (nios2_2nd_core_custom_instruction_master_multi_readrb),                         //                .multi_readrb
		.ci_slave_multi_writerc    (nios2_2nd_core_custom_instruction_master_multi_writerc),                        //                .multi_writerc
		.ci_slave_multi_a          (nios2_2nd_core_custom_instruction_master_multi_a),                              //                .multi_a
		.ci_slave_multi_b          (nios2_2nd_core_custom_instruction_master_multi_b),                              //                .multi_b
		.ci_slave_multi_c          (nios2_2nd_core_custom_instruction_master_multi_c),                              //                .multi_c
		.comb_ci_master_result     (),                                                                              //  comb_ci_master.result
		.multi_ci_master_clk       (nios2_2nd_core_custom_instruction_master_translator_multi_ci_master_clk),       // multi_ci_master.clk
		.multi_ci_master_reset     (nios2_2nd_core_custom_instruction_master_translator_multi_ci_master_reset),     //                .reset
		.multi_ci_master_clken     (nios2_2nd_core_custom_instruction_master_translator_multi_ci_master_clk_en),    //                .clk_en
		.multi_ci_master_reset_req (nios2_2nd_core_custom_instruction_master_translator_multi_ci_master_reset_req), //                .reset_req
		.multi_ci_master_start     (nios2_2nd_core_custom_instruction_master_translator_multi_ci_master_start),     //                .start
		.multi_ci_master_done      (nios2_2nd_core_custom_instruction_master_translator_multi_ci_master_done),      //                .done
		.multi_ci_master_dataa     (nios2_2nd_core_custom_instruction_master_translator_multi_ci_master_dataa),     //                .dataa
		.multi_ci_master_datab     (nios2_2nd_core_custom_instruction_master_translator_multi_ci_master_datab),     //                .datab
		.multi_ci_master_result    (nios2_2nd_core_custom_instruction_master_translator_multi_ci_master_result),    //                .result
		.multi_ci_master_n         (nios2_2nd_core_custom_instruction_master_translator_multi_ci_master_n),         //                .n
		.multi_ci_master_readra    (nios2_2nd_core_custom_instruction_master_translator_multi_ci_master_readra),    //                .readra
		.multi_ci_master_readrb    (nios2_2nd_core_custom_instruction_master_translator_multi_ci_master_readrb),    //                .readrb
		.multi_ci_master_writerc   (nios2_2nd_core_custom_instruction_master_translator_multi_ci_master_writerc),   //                .writerc
		.multi_ci_master_a         (nios2_2nd_core_custom_instruction_master_translator_multi_ci_master_a),         //                .a
		.multi_ci_master_b         (nios2_2nd_core_custom_instruction_master_translator_multi_ci_master_b),         //                .b
		.multi_ci_master_c         (nios2_2nd_core_custom_instruction_master_translator_multi_ci_master_c),         //                .c
		.ci_slave_dataa            (32'b00000000000000000000000000000000),                                          //     (terminated)
		.ci_slave_datab            (32'b00000000000000000000000000000000),                                          //     (terminated)
		.ci_slave_n                (8'b00000000),                                                                   //     (terminated)
		.ci_slave_readra           (1'b0),                                                                          //     (terminated)
		.ci_slave_readrb           (1'b0),                                                                          //     (terminated)
		.ci_slave_writerc          (1'b0),                                                                          //     (terminated)
		.ci_slave_a                (5'b00000),                                                                      //     (terminated)
		.ci_slave_b                (5'b00000),                                                                      //     (terminated)
		.ci_slave_c                (5'b00000),                                                                      //     (terminated)
		.ci_slave_ipending         (32'b00000000000000000000000000000000),                                          //     (terminated)
		.ci_slave_estatus          (1'b0),                                                                          //     (terminated)
		.comb_ci_master_dataa      (),                                                                              //     (terminated)
		.comb_ci_master_datab      (),                                                                              //     (terminated)
		.comb_ci_master_n          (),                                                                              //     (terminated)
		.comb_ci_master_readra     (),                                                                              //     (terminated)
		.comb_ci_master_readrb     (),                                                                              //     (terminated)
		.comb_ci_master_writerc    (),                                                                              //     (terminated)
		.comb_ci_master_a          (),                                                                              //     (terminated)
		.comb_ci_master_b          (),                                                                              //     (terminated)
		.comb_ci_master_c          (),                                                                              //     (terminated)
		.comb_ci_master_ipending   (),                                                                              //     (terminated)
		.comb_ci_master_estatus    ()                                                                               //     (terminated)
	);

	Computer_System_Nios2_2nd_Core_custom_instruction_master_multi_xconnect nios2_2nd_core_custom_instruction_master_multi_xconnect (
		.ci_slave_dataa       (nios2_2nd_core_custom_instruction_master_translator_multi_ci_master_dataa),     //   ci_slave.dataa
		.ci_slave_datab       (nios2_2nd_core_custom_instruction_master_translator_multi_ci_master_datab),     //           .datab
		.ci_slave_result      (nios2_2nd_core_custom_instruction_master_translator_multi_ci_master_result),    //           .result
		.ci_slave_n           (nios2_2nd_core_custom_instruction_master_translator_multi_ci_master_n),         //           .n
		.ci_slave_readra      (nios2_2nd_core_custom_instruction_master_translator_multi_ci_master_readra),    //           .readra
		.ci_slave_readrb      (nios2_2nd_core_custom_instruction_master_translator_multi_ci_master_readrb),    //           .readrb
		.ci_slave_writerc     (nios2_2nd_core_custom_instruction_master_translator_multi_ci_master_writerc),   //           .writerc
		.ci_slave_a           (nios2_2nd_core_custom_instruction_master_translator_multi_ci_master_a),         //           .a
		.ci_slave_b           (nios2_2nd_core_custom_instruction_master_translator_multi_ci_master_b),         //           .b
		.ci_slave_c           (nios2_2nd_core_custom_instruction_master_translator_multi_ci_master_c),         //           .c
		.ci_slave_ipending    (),                                                                              //           .ipending
		.ci_slave_estatus     (),                                                                              //           .estatus
		.ci_slave_clk         (nios2_2nd_core_custom_instruction_master_translator_multi_ci_master_clk),       //           .clk
		.ci_slave_reset       (nios2_2nd_core_custom_instruction_master_translator_multi_ci_master_reset),     //           .reset
		.ci_slave_clken       (nios2_2nd_core_custom_instruction_master_translator_multi_ci_master_clk_en),    //           .clk_en
		.ci_slave_reset_req   (nios2_2nd_core_custom_instruction_master_translator_multi_ci_master_reset_req), //           .reset_req
		.ci_slave_start       (nios2_2nd_core_custom_instruction_master_translator_multi_ci_master_start),     //           .start
		.ci_slave_done        (nios2_2nd_core_custom_instruction_master_translator_multi_ci_master_done),      //           .done
		.ci_master0_dataa     (nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_dataa),      // ci_master0.dataa
		.ci_master0_datab     (nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_datab),      //           .datab
		.ci_master0_result    (nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_result),     //           .result
		.ci_master0_n         (nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_n),          //           .n
		.ci_master0_readra    (nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_readra),     //           .readra
		.ci_master0_readrb    (nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_readrb),     //           .readrb
		.ci_master0_writerc   (nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_writerc),    //           .writerc
		.ci_master0_a         (nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_a),          //           .a
		.ci_master0_b         (nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_b),          //           .b
		.ci_master0_c         (nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_c),          //           .c
		.ci_master0_ipending  (nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_ipending),   //           .ipending
		.ci_master0_estatus   (nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_estatus),    //           .estatus
		.ci_master0_clk       (nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_clk),        //           .clk
		.ci_master0_reset     (nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_reset),      //           .reset
		.ci_master0_clken     (nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_clk_en),     //           .clk_en
		.ci_master0_reset_req (nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_reset_req),  //           .reset_req
		.ci_master0_start     (nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_start),      //           .start
		.ci_master0_done      (nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_done)        //           .done
	);

	altera_customins_slave_translator #(
		.N_WIDTH          (2),
		.USE_DONE         (1),
		.NUM_FIXED_CYCLES (1)
	) nios2_2nd_core_custom_instruction_master_multi_slave_translator0 (
		.ci_slave_dataa      (nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_dataa),          //  ci_slave.dataa
		.ci_slave_datab      (nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_datab),          //          .datab
		.ci_slave_result     (nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_result),         //          .result
		.ci_slave_n          (nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_n),              //          .n
		.ci_slave_readra     (nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_readra),         //          .readra
		.ci_slave_readrb     (nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_readrb),         //          .readrb
		.ci_slave_writerc    (nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_writerc),        //          .writerc
		.ci_slave_a          (nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_a),              //          .a
		.ci_slave_b          (nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_b),              //          .b
		.ci_slave_c          (nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_c),              //          .c
		.ci_slave_ipending   (nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_ipending),       //          .ipending
		.ci_slave_estatus    (nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_estatus),        //          .estatus
		.ci_slave_clk        (nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_clk),            //          .clk
		.ci_slave_clken      (nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_clk_en),         //          .clk_en
		.ci_slave_reset_req  (nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_reset_req),      //          .reset_req
		.ci_slave_reset      (nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_reset),          //          .reset
		.ci_slave_start      (nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_start),          //          .start
		.ci_slave_done       (nios2_2nd_core_custom_instruction_master_multi_xconnect_ci_master0_done),           //          .done
		.ci_master_dataa     (nios2_2nd_core_custom_instruction_master_multi_slave_translator0_ci_master_dataa),  // ci_master.dataa
		.ci_master_datab     (nios2_2nd_core_custom_instruction_master_multi_slave_translator0_ci_master_datab),  //          .datab
		.ci_master_result    (nios2_2nd_core_custom_instruction_master_multi_slave_translator0_ci_master_result), //          .result
		.ci_master_n         (nios2_2nd_core_custom_instruction_master_multi_slave_translator0_ci_master_n),      //          .n
		.ci_master_clk       (nios2_2nd_core_custom_instruction_master_multi_slave_translator0_ci_master_clk),    //          .clk
		.ci_master_clken     (nios2_2nd_core_custom_instruction_master_multi_slave_translator0_ci_master_clk_en), //          .clk_en
		.ci_master_reset     (nios2_2nd_core_custom_instruction_master_multi_slave_translator0_ci_master_reset),  //          .reset
		.ci_master_start     (nios2_2nd_core_custom_instruction_master_multi_slave_translator0_ci_master_start),  //          .start
		.ci_master_done      (nios2_2nd_core_custom_instruction_master_multi_slave_translator0_ci_master_done),   //          .done
		.ci_master_readra    (),                                                                                  // (terminated)
		.ci_master_readrb    (),                                                                                  // (terminated)
		.ci_master_writerc   (),                                                                                  // (terminated)
		.ci_master_a         (),                                                                                  // (terminated)
		.ci_master_b         (),                                                                                  // (terminated)
		.ci_master_c         (),                                                                                  // (terminated)
		.ci_master_ipending  (),                                                                                  // (terminated)
		.ci_master_estatus   (),                                                                                  // (terminated)
		.ci_master_reset_req ()                                                                                   // (terminated)
	);

	Computer_System_mm_interconnect_0 mm_interconnect_0 (
		.System_PLL_sys_clk_clk                                              (system_pll_sys_clk_clk),                                                                //                                       System_PLL_sys_clk.clk
		.AV_Config_reset_reset_bridge_in_reset_reset                         (rst_controller_reset_out_reset),                                                        //                    AV_Config_reset_reset_bridge_in_reset.reset
		.JTAG_to_FPGA_Bridge_clk_reset_reset_bridge_in_reset_reset           (rst_controller_reset_out_reset),                                                        //      JTAG_to_FPGA_Bridge_clk_reset_reset_bridge_in_reset.reset
		.Nios2_2nd_Core_reset_reset_bridge_in_reset_reset                    (rst_controller_002_reset_out_reset),                                                    //               Nios2_2nd_Core_reset_reset_bridge_in_reset.reset
		.Nios2_reset_reset_bridge_in_reset_reset                             (rst_controller_001_reset_out_reset),                                                    //                        Nios2_reset_reset_bridge_in_reset.reset
		.JTAG_to_FPGA_Bridge_master_address                                  (jtag_to_fpga_bridge_master_address),                                                    //                               JTAG_to_FPGA_Bridge_master.address
		.JTAG_to_FPGA_Bridge_master_waitrequest                              (jtag_to_fpga_bridge_master_waitrequest),                                                //                                                         .waitrequest
		.JTAG_to_FPGA_Bridge_master_byteenable                               (jtag_to_fpga_bridge_master_byteenable),                                                 //                                                         .byteenable
		.JTAG_to_FPGA_Bridge_master_read                                     (jtag_to_fpga_bridge_master_read),                                                       //                                                         .read
		.JTAG_to_FPGA_Bridge_master_readdata                                 (jtag_to_fpga_bridge_master_readdata),                                                   //                                                         .readdata
		.JTAG_to_FPGA_Bridge_master_readdatavalid                            (jtag_to_fpga_bridge_master_readdatavalid),                                              //                                                         .readdatavalid
		.JTAG_to_FPGA_Bridge_master_write                                    (jtag_to_fpga_bridge_master_write),                                                      //                                                         .write
		.JTAG_to_FPGA_Bridge_master_writedata                                (jtag_to_fpga_bridge_master_writedata),                                                  //                                                         .writedata
		.Nios2_data_master_address                                           (nios2_data_master_address),                                                             //                                        Nios2_data_master.address
		.Nios2_data_master_waitrequest                                       (nios2_data_master_waitrequest),                                                         //                                                         .waitrequest
		.Nios2_data_master_byteenable                                        (nios2_data_master_byteenable),                                                          //                                                         .byteenable
		.Nios2_data_master_read                                              (nios2_data_master_read),                                                                //                                                         .read
		.Nios2_data_master_readdata                                          (nios2_data_master_readdata),                                                            //                                                         .readdata
		.Nios2_data_master_write                                             (nios2_data_master_write),                                                               //                                                         .write
		.Nios2_data_master_writedata                                         (nios2_data_master_writedata),                                                           //                                                         .writedata
		.Nios2_data_master_debugaccess                                       (nios2_data_master_debugaccess),                                                         //                                                         .debugaccess
		.Nios2_instruction_master_address                                    (nios2_instruction_master_address),                                                      //                                 Nios2_instruction_master.address
		.Nios2_instruction_master_waitrequest                                (nios2_instruction_master_waitrequest),                                                  //                                                         .waitrequest
		.Nios2_instruction_master_read                                       (nios2_instruction_master_read),                                                         //                                                         .read
		.Nios2_instruction_master_readdata                                   (nios2_instruction_master_readdata),                                                     //                                                         .readdata
		.Nios2_instruction_master_readdatavalid                              (nios2_instruction_master_readdatavalid),                                                //                                                         .readdatavalid
		.Nios2_2nd_Core_data_master_address                                  (nios2_2nd_core_data_master_address),                                                    //                               Nios2_2nd_Core_data_master.address
		.Nios2_2nd_Core_data_master_waitrequest                              (nios2_2nd_core_data_master_waitrequest),                                                //                                                         .waitrequest
		.Nios2_2nd_Core_data_master_byteenable                               (nios2_2nd_core_data_master_byteenable),                                                 //                                                         .byteenable
		.Nios2_2nd_Core_data_master_read                                     (nios2_2nd_core_data_master_read),                                                       //                                                         .read
		.Nios2_2nd_Core_data_master_readdata                                 (nios2_2nd_core_data_master_readdata),                                                   //                                                         .readdata
		.Nios2_2nd_Core_data_master_write                                    (nios2_2nd_core_data_master_write),                                                      //                                                         .write
		.Nios2_2nd_Core_data_master_writedata                                (nios2_2nd_core_data_master_writedata),                                                  //                                                         .writedata
		.Nios2_2nd_Core_data_master_debugaccess                              (nios2_2nd_core_data_master_debugaccess),                                                //                                                         .debugaccess
		.Nios2_2nd_Core_instruction_master_address                           (nios2_2nd_core_instruction_master_address),                                             //                        Nios2_2nd_Core_instruction_master.address
		.Nios2_2nd_Core_instruction_master_waitrequest                       (nios2_2nd_core_instruction_master_waitrequest),                                         //                                                         .waitrequest
		.Nios2_2nd_Core_instruction_master_read                              (nios2_2nd_core_instruction_master_read),                                                //                                                         .read
		.Nios2_2nd_Core_instruction_master_readdata                          (nios2_2nd_core_instruction_master_readdata),                                            //                                                         .readdata
		.Nios2_2nd_Core_instruction_master_readdatavalid                     (nios2_2nd_core_instruction_master_readdatavalid),                                       //                                                         .readdatavalid
		.VGA_Subsystem_pixel_dma_master_address                              (vga_subsystem_pixel_dma_master_address),                                                //                           VGA_Subsystem_pixel_dma_master.address
		.VGA_Subsystem_pixel_dma_master_waitrequest                          (vga_subsystem_pixel_dma_master_waitrequest),                                            //                                                         .waitrequest
		.VGA_Subsystem_pixel_dma_master_read                                 (vga_subsystem_pixel_dma_master_read),                                                   //                                                         .read
		.VGA_Subsystem_pixel_dma_master_readdata                             (vga_subsystem_pixel_dma_master_readdata),                                               //                                                         .readdata
		.VGA_Subsystem_pixel_dma_master_readdatavalid                        (vga_subsystem_pixel_dma_master_readdatavalid),                                          //                                                         .readdatavalid
		.VGA_Subsystem_pixel_dma_master_lock                                 (vga_subsystem_pixel_dma_master_lock),                                                   //                                                         .lock
		.Video_In_Subsystem_video_in_dma_master_address                      (video_in_subsystem_video_in_dma_master_address),                                        //                   Video_In_Subsystem_video_in_dma_master.address
		.Video_In_Subsystem_video_in_dma_master_waitrequest                  (video_in_subsystem_video_in_dma_master_waitrequest),                                    //                                                         .waitrequest
		.Video_In_Subsystem_video_in_dma_master_write                        (video_in_subsystem_video_in_dma_master_write),                                          //                                                         .write
		.Video_In_Subsystem_video_in_dma_master_writedata                    (video_in_subsystem_video_in_dma_master_writedata),                                      //                                                         .writedata
		.Audio_Subsystem_audio_slave_address                                 (mm_interconnect_0_audio_subsystem_audio_slave_address),                                 //                              Audio_Subsystem_audio_slave.address
		.Audio_Subsystem_audio_slave_write                                   (mm_interconnect_0_audio_subsystem_audio_slave_write),                                   //                                                         .write
		.Audio_Subsystem_audio_slave_read                                    (mm_interconnect_0_audio_subsystem_audio_slave_read),                                    //                                                         .read
		.Audio_Subsystem_audio_slave_readdata                                (mm_interconnect_0_audio_subsystem_audio_slave_readdata),                                //                                                         .readdata
		.Audio_Subsystem_audio_slave_writedata                               (mm_interconnect_0_audio_subsystem_audio_slave_writedata),                               //                                                         .writedata
		.Audio_Subsystem_audio_slave_chipselect                              (mm_interconnect_0_audio_subsystem_audio_slave_chipselect),                              //                                                         .chipselect
		.AV_Config_avalon_av_config_slave_address                            (mm_interconnect_0_av_config_avalon_av_config_slave_address),                            //                         AV_Config_avalon_av_config_slave.address
		.AV_Config_avalon_av_config_slave_write                              (mm_interconnect_0_av_config_avalon_av_config_slave_write),                              //                                                         .write
		.AV_Config_avalon_av_config_slave_read                               (mm_interconnect_0_av_config_avalon_av_config_slave_read),                               //                                                         .read
		.AV_Config_avalon_av_config_slave_readdata                           (mm_interconnect_0_av_config_avalon_av_config_slave_readdata),                           //                                                         .readdata
		.AV_Config_avalon_av_config_slave_writedata                          (mm_interconnect_0_av_config_avalon_av_config_slave_writedata),                          //                                                         .writedata
		.AV_Config_avalon_av_config_slave_byteenable                         (mm_interconnect_0_av_config_avalon_av_config_slave_byteenable),                         //                                                         .byteenable
		.AV_Config_avalon_av_config_slave_waitrequest                        (mm_interconnect_0_av_config_avalon_av_config_slave_waitrequest),                        //                                                         .waitrequest
		.Char_LCD_16x2_avalon_lcd_slave_address                              (mm_interconnect_0_char_lcd_16x2_avalon_lcd_slave_address),                              //                           Char_LCD_16x2_avalon_lcd_slave.address
		.Char_LCD_16x2_avalon_lcd_slave_write                                (mm_interconnect_0_char_lcd_16x2_avalon_lcd_slave_write),                                //                                                         .write
		.Char_LCD_16x2_avalon_lcd_slave_read                                 (mm_interconnect_0_char_lcd_16x2_avalon_lcd_slave_read),                                 //                                                         .read
		.Char_LCD_16x2_avalon_lcd_slave_readdata                             (mm_interconnect_0_char_lcd_16x2_avalon_lcd_slave_readdata),                             //                                                         .readdata
		.Char_LCD_16x2_avalon_lcd_slave_writedata                            (mm_interconnect_0_char_lcd_16x2_avalon_lcd_slave_writedata),                            //                                                         .writedata
		.Char_LCD_16x2_avalon_lcd_slave_waitrequest                          (mm_interconnect_0_char_lcd_16x2_avalon_lcd_slave_waitrequest),                          //                                                         .waitrequest
		.Char_LCD_16x2_avalon_lcd_slave_chipselect                           (mm_interconnect_0_char_lcd_16x2_avalon_lcd_slave_chipselect),                           //                                                         .chipselect
		.Expansion_JP5_s1_address                                            (mm_interconnect_0_expansion_jp5_s1_address),                                            //                                         Expansion_JP5_s1.address
		.Expansion_JP5_s1_write                                              (mm_interconnect_0_expansion_jp5_s1_write),                                              //                                                         .write
		.Expansion_JP5_s1_readdata                                           (mm_interconnect_0_expansion_jp5_s1_readdata),                                           //                                                         .readdata
		.Expansion_JP5_s1_writedata                                          (mm_interconnect_0_expansion_jp5_s1_writedata),                                          //                                                         .writedata
		.Expansion_JP5_s1_chipselect                                         (mm_interconnect_0_expansion_jp5_s1_chipselect),                                         //                                                         .chipselect
		.Flash_flash_data_address                                            (mm_interconnect_0_flash_flash_data_address),                                            //                                         Flash_flash_data.address
		.Flash_flash_data_write                                              (mm_interconnect_0_flash_flash_data_write),                                              //                                                         .write
		.Flash_flash_data_read                                               (mm_interconnect_0_flash_flash_data_read),                                               //                                                         .read
		.Flash_flash_data_readdata                                           (mm_interconnect_0_flash_flash_data_readdata),                                           //                                                         .readdata
		.Flash_flash_data_writedata                                          (mm_interconnect_0_flash_flash_data_writedata),                                          //                                                         .writedata
		.Flash_flash_data_byteenable                                         (mm_interconnect_0_flash_flash_data_byteenable),                                         //                                                         .byteenable
		.Flash_flash_data_waitrequest                                        (mm_interconnect_0_flash_flash_data_waitrequest),                                        //                                                         .waitrequest
		.Flash_flash_data_chipselect                                         (mm_interconnect_0_flash_flash_data_chipselect),                                         //                                                         .chipselect
		.Flash_flash_erase_control_write                                     (mm_interconnect_0_flash_flash_erase_control_write),                                     //                                Flash_flash_erase_control.write
		.Flash_flash_erase_control_read                                      (mm_interconnect_0_flash_flash_erase_control_read),                                      //                                                         .read
		.Flash_flash_erase_control_readdata                                  (mm_interconnect_0_flash_flash_erase_control_readdata),                                  //                                                         .readdata
		.Flash_flash_erase_control_writedata                                 (mm_interconnect_0_flash_flash_erase_control_writedata),                                 //                                                         .writedata
		.Flash_flash_erase_control_byteenable                                (mm_interconnect_0_flash_flash_erase_control_byteenable),                                //                                                         .byteenable
		.Flash_flash_erase_control_waitrequest                               (mm_interconnect_0_flash_flash_erase_control_waitrequest),                               //                                                         .waitrequest
		.Flash_flash_erase_control_chipselect                                (mm_interconnect_0_flash_flash_erase_control_chipselect),                                //                                                         .chipselect
		.Green_LEDs_s1_address                                               (mm_interconnect_0_green_leds_s1_address),                                               //                                            Green_LEDs_s1.address
		.Green_LEDs_s1_write                                                 (mm_interconnect_0_green_leds_s1_write),                                                 //                                                         .write
		.Green_LEDs_s1_readdata                                              (mm_interconnect_0_green_leds_s1_readdata),                                              //                                                         .readdata
		.Green_LEDs_s1_writedata                                             (mm_interconnect_0_green_leds_s1_writedata),                                             //                                                         .writedata
		.Green_LEDs_s1_chipselect                                            (mm_interconnect_0_green_leds_s1_chipselect),                                            //                                                         .chipselect
		.HEX3_HEX0_s1_address                                                (mm_interconnect_0_hex3_hex0_s1_address),                                                //                                             HEX3_HEX0_s1.address
		.HEX3_HEX0_s1_write                                                  (mm_interconnect_0_hex3_hex0_s1_write),                                                  //                                                         .write
		.HEX3_HEX0_s1_readdata                                               (mm_interconnect_0_hex3_hex0_s1_readdata),                                               //                                                         .readdata
		.HEX3_HEX0_s1_writedata                                              (mm_interconnect_0_hex3_hex0_s1_writedata),                                              //                                                         .writedata
		.HEX3_HEX0_s1_chipselect                                             (mm_interconnect_0_hex3_hex0_s1_chipselect),                                             //                                                         .chipselect
		.HEX7_HEX4_s1_address                                                (mm_interconnect_0_hex7_hex4_s1_address),                                                //                                             HEX7_HEX4_s1.address
		.HEX7_HEX4_s1_write                                                  (mm_interconnect_0_hex7_hex4_s1_write),                                                  //                                                         .write
		.HEX7_HEX4_s1_readdata                                               (mm_interconnect_0_hex7_hex4_s1_readdata),                                               //                                                         .readdata
		.HEX7_HEX4_s1_writedata                                              (mm_interconnect_0_hex7_hex4_s1_writedata),                                              //                                                         .writedata
		.HEX7_HEX4_s1_chipselect                                             (mm_interconnect_0_hex7_hex4_s1_chipselect),                                             //                                                         .chipselect
		.Interval_Timer_s1_address                                           (mm_interconnect_0_interval_timer_s1_address),                                           //                                        Interval_Timer_s1.address
		.Interval_Timer_s1_write                                             (mm_interconnect_0_interval_timer_s1_write),                                             //                                                         .write
		.Interval_Timer_s1_readdata                                          (mm_interconnect_0_interval_timer_s1_readdata),                                          //                                                         .readdata
		.Interval_Timer_s1_writedata                                         (mm_interconnect_0_interval_timer_s1_writedata),                                         //                                                         .writedata
		.Interval_Timer_s1_chipselect                                        (mm_interconnect_0_interval_timer_s1_chipselect),                                        //                                                         .chipselect
		.Interval_Timer_2_s1_address                                         (mm_interconnect_0_interval_timer_2_s1_address),                                         //                                      Interval_Timer_2_s1.address
		.Interval_Timer_2_s1_write                                           (mm_interconnect_0_interval_timer_2_s1_write),                                           //                                                         .write
		.Interval_Timer_2_s1_readdata                                        (mm_interconnect_0_interval_timer_2_s1_readdata),                                        //                                                         .readdata
		.Interval_Timer_2_s1_writedata                                       (mm_interconnect_0_interval_timer_2_s1_writedata),                                       //                                                         .writedata
		.Interval_Timer_2_s1_chipselect                                      (mm_interconnect_0_interval_timer_2_s1_chipselect),                                      //                                                         .chipselect
		.Interval_Timer_2nd_Core_s1_address                                  (mm_interconnect_0_interval_timer_2nd_core_s1_address),                                  //                               Interval_Timer_2nd_Core_s1.address
		.Interval_Timer_2nd_Core_s1_write                                    (mm_interconnect_0_interval_timer_2nd_core_s1_write),                                    //                                                         .write
		.Interval_Timer_2nd_Core_s1_readdata                                 (mm_interconnect_0_interval_timer_2nd_core_s1_readdata),                                 //                                                         .readdata
		.Interval_Timer_2nd_Core_s1_writedata                                (mm_interconnect_0_interval_timer_2nd_core_s1_writedata),                                //                                                         .writedata
		.Interval_Timer_2nd_Core_s1_chipselect                               (mm_interconnect_0_interval_timer_2nd_core_s1_chipselect),                               //                                                         .chipselect
		.Interval_Timer_2nd_Core_2_s1_address                                (mm_interconnect_0_interval_timer_2nd_core_2_s1_address),                                //                             Interval_Timer_2nd_Core_2_s1.address
		.Interval_Timer_2nd_Core_2_s1_write                                  (mm_interconnect_0_interval_timer_2nd_core_2_s1_write),                                  //                                                         .write
		.Interval_Timer_2nd_Core_2_s1_readdata                               (mm_interconnect_0_interval_timer_2nd_core_2_s1_readdata),                               //                                                         .readdata
		.Interval_Timer_2nd_Core_2_s1_writedata                              (mm_interconnect_0_interval_timer_2nd_core_2_s1_writedata),                              //                                                         .writedata
		.Interval_Timer_2nd_Core_2_s1_chipselect                             (mm_interconnect_0_interval_timer_2nd_core_2_s1_chipselect),                             //                                                         .chipselect
		.IrDA_avalon_irda_slave_address                                      (mm_interconnect_0_irda_avalon_irda_slave_address),                                      //                                   IrDA_avalon_irda_slave.address
		.IrDA_avalon_irda_slave_write                                        (mm_interconnect_0_irda_avalon_irda_slave_write),                                        //                                                         .write
		.IrDA_avalon_irda_slave_read                                         (mm_interconnect_0_irda_avalon_irda_slave_read),                                         //                                                         .read
		.IrDA_avalon_irda_slave_readdata                                     (mm_interconnect_0_irda_avalon_irda_slave_readdata),                                     //                                                         .readdata
		.IrDA_avalon_irda_slave_writedata                                    (mm_interconnect_0_irda_avalon_irda_slave_writedata),                                    //                                                         .writedata
		.IrDA_avalon_irda_slave_byteenable                                   (mm_interconnect_0_irda_avalon_irda_slave_byteenable),                                   //                                                         .byteenable
		.IrDA_avalon_irda_slave_chipselect                                   (mm_interconnect_0_irda_avalon_irda_slave_chipselect),                                   //                                                         .chipselect
		.JTAG_UART_avalon_jtag_slave_address                                 (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),                                 //                              JTAG_UART_avalon_jtag_slave.address
		.JTAG_UART_avalon_jtag_slave_write                                   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),                                   //                                                         .write
		.JTAG_UART_avalon_jtag_slave_read                                    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),                                    //                                                         .read
		.JTAG_UART_avalon_jtag_slave_readdata                                (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),                                //                                                         .readdata
		.JTAG_UART_avalon_jtag_slave_writedata                               (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),                               //                                                         .writedata
		.JTAG_UART_avalon_jtag_slave_waitrequest                             (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest),                             //                                                         .waitrequest
		.JTAG_UART_avalon_jtag_slave_chipselect                              (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),                              //                                                         .chipselect
		.JTAG_UART_2nd_Core_avalon_jtag_slave_address                        (mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_address),                        //                     JTAG_UART_2nd_Core_avalon_jtag_slave.address
		.JTAG_UART_2nd_Core_avalon_jtag_slave_write                          (mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_write),                          //                                                         .write
		.JTAG_UART_2nd_Core_avalon_jtag_slave_read                           (mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_read),                           //                                                         .read
		.JTAG_UART_2nd_Core_avalon_jtag_slave_readdata                       (mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_readdata),                       //                                                         .readdata
		.JTAG_UART_2nd_Core_avalon_jtag_slave_writedata                      (mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_writedata),                      //                                                         .writedata
		.JTAG_UART_2nd_Core_avalon_jtag_slave_waitrequest                    (mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_waitrequest),                    //                                                         .waitrequest
		.JTAG_UART_2nd_Core_avalon_jtag_slave_chipselect                     (mm_interconnect_0_jtag_uart_2nd_core_avalon_jtag_slave_chipselect),                     //                                                         .chipselect
		.Nios2_debug_mem_slave_address                                       (mm_interconnect_0_nios2_debug_mem_slave_address),                                       //                                    Nios2_debug_mem_slave.address
		.Nios2_debug_mem_slave_write                                         (mm_interconnect_0_nios2_debug_mem_slave_write),                                         //                                                         .write
		.Nios2_debug_mem_slave_read                                          (mm_interconnect_0_nios2_debug_mem_slave_read),                                          //                                                         .read
		.Nios2_debug_mem_slave_readdata                                      (mm_interconnect_0_nios2_debug_mem_slave_readdata),                                      //                                                         .readdata
		.Nios2_debug_mem_slave_writedata                                     (mm_interconnect_0_nios2_debug_mem_slave_writedata),                                     //                                                         .writedata
		.Nios2_debug_mem_slave_byteenable                                    (mm_interconnect_0_nios2_debug_mem_slave_byteenable),                                    //                                                         .byteenable
		.Nios2_debug_mem_slave_waitrequest                                   (mm_interconnect_0_nios2_debug_mem_slave_waitrequest),                                   //                                                         .waitrequest
		.Nios2_debug_mem_slave_debugaccess                                   (mm_interconnect_0_nios2_debug_mem_slave_debugaccess),                                   //                                                         .debugaccess
		.Nios2_2nd_Core_debug_mem_slave_address                              (mm_interconnect_0_nios2_2nd_core_debug_mem_slave_address),                              //                           Nios2_2nd_Core_debug_mem_slave.address
		.Nios2_2nd_Core_debug_mem_slave_write                                (mm_interconnect_0_nios2_2nd_core_debug_mem_slave_write),                                //                                                         .write
		.Nios2_2nd_Core_debug_mem_slave_read                                 (mm_interconnect_0_nios2_2nd_core_debug_mem_slave_read),                                 //                                                         .read
		.Nios2_2nd_Core_debug_mem_slave_readdata                             (mm_interconnect_0_nios2_2nd_core_debug_mem_slave_readdata),                             //                                                         .readdata
		.Nios2_2nd_Core_debug_mem_slave_writedata                            (mm_interconnect_0_nios2_2nd_core_debug_mem_slave_writedata),                            //                                                         .writedata
		.Nios2_2nd_Core_debug_mem_slave_byteenable                           (mm_interconnect_0_nios2_2nd_core_debug_mem_slave_byteenable),                           //                                                         .byteenable
		.Nios2_2nd_Core_debug_mem_slave_waitrequest                          (mm_interconnect_0_nios2_2nd_core_debug_mem_slave_waitrequest),                          //                                                         .waitrequest
		.Nios2_2nd_Core_debug_mem_slave_debugaccess                          (mm_interconnect_0_nios2_2nd_core_debug_mem_slave_debugaccess),                          //                                                         .debugaccess
		.PS2_Port_avalon_ps2_slave_address                                   (mm_interconnect_0_ps2_port_avalon_ps2_slave_address),                                   //                                PS2_Port_avalon_ps2_slave.address
		.PS2_Port_avalon_ps2_slave_write                                     (mm_interconnect_0_ps2_port_avalon_ps2_slave_write),                                     //                                                         .write
		.PS2_Port_avalon_ps2_slave_read                                      (mm_interconnect_0_ps2_port_avalon_ps2_slave_read),                                      //                                                         .read
		.PS2_Port_avalon_ps2_slave_readdata                                  (mm_interconnect_0_ps2_port_avalon_ps2_slave_readdata),                                  //                                                         .readdata
		.PS2_Port_avalon_ps2_slave_writedata                                 (mm_interconnect_0_ps2_port_avalon_ps2_slave_writedata),                                 //                                                         .writedata
		.PS2_Port_avalon_ps2_slave_byteenable                                (mm_interconnect_0_ps2_port_avalon_ps2_slave_byteenable),                                //                                                         .byteenable
		.PS2_Port_avalon_ps2_slave_waitrequest                               (mm_interconnect_0_ps2_port_avalon_ps2_slave_waitrequest),                               //                                                         .waitrequest
		.PS2_Port_avalon_ps2_slave_chipselect                                (mm_interconnect_0_ps2_port_avalon_ps2_slave_chipselect),                                //                                                         .chipselect
		.PS2_Port_Dual_avalon_ps2_slave_address                              (mm_interconnect_0_ps2_port_dual_avalon_ps2_slave_address),                              //                           PS2_Port_Dual_avalon_ps2_slave.address
		.PS2_Port_Dual_avalon_ps2_slave_write                                (mm_interconnect_0_ps2_port_dual_avalon_ps2_slave_write),                                //                                                         .write
		.PS2_Port_Dual_avalon_ps2_slave_read                                 (mm_interconnect_0_ps2_port_dual_avalon_ps2_slave_read),                                 //                                                         .read
		.PS2_Port_Dual_avalon_ps2_slave_readdata                             (mm_interconnect_0_ps2_port_dual_avalon_ps2_slave_readdata),                             //                                                         .readdata
		.PS2_Port_Dual_avalon_ps2_slave_writedata                            (mm_interconnect_0_ps2_port_dual_avalon_ps2_slave_writedata),                            //                                                         .writedata
		.PS2_Port_Dual_avalon_ps2_slave_byteenable                           (mm_interconnect_0_ps2_port_dual_avalon_ps2_slave_byteenable),                           //                                                         .byteenable
		.PS2_Port_Dual_avalon_ps2_slave_waitrequest                          (mm_interconnect_0_ps2_port_dual_avalon_ps2_slave_waitrequest),                          //                                                         .waitrequest
		.PS2_Port_Dual_avalon_ps2_slave_chipselect                           (mm_interconnect_0_ps2_port_dual_avalon_ps2_slave_chipselect),                           //                                                         .chipselect
		.Pushbuttons_s1_address                                              (mm_interconnect_0_pushbuttons_s1_address),                                              //                                           Pushbuttons_s1.address
		.Pushbuttons_s1_write                                                (mm_interconnect_0_pushbuttons_s1_write),                                                //                                                         .write
		.Pushbuttons_s1_readdata                                             (mm_interconnect_0_pushbuttons_s1_readdata),                                             //                                                         .readdata
		.Pushbuttons_s1_writedata                                            (mm_interconnect_0_pushbuttons_s1_writedata),                                            //                                                         .writedata
		.Pushbuttons_s1_chipselect                                           (mm_interconnect_0_pushbuttons_s1_chipselect),                                           //                                                         .chipselect
		.Red_LEDs_s1_address                                                 (mm_interconnect_0_red_leds_s1_address),                                                 //                                              Red_LEDs_s1.address
		.Red_LEDs_s1_write                                                   (mm_interconnect_0_red_leds_s1_write),                                                   //                                                         .write
		.Red_LEDs_s1_readdata                                                (mm_interconnect_0_red_leds_s1_readdata),                                                //                                                         .readdata
		.Red_LEDs_s1_writedata                                               (mm_interconnect_0_red_leds_s1_writedata),                                               //                                                         .writedata
		.Red_LEDs_s1_chipselect                                              (mm_interconnect_0_red_leds_s1_chipselect),                                              //                                                         .chipselect
		.SD_Card_avalon_sdcard_slave_address                                 (mm_interconnect_0_sd_card_avalon_sdcard_slave_address),                                 //                              SD_Card_avalon_sdcard_slave.address
		.SD_Card_avalon_sdcard_slave_write                                   (mm_interconnect_0_sd_card_avalon_sdcard_slave_write),                                   //                                                         .write
		.SD_Card_avalon_sdcard_slave_read                                    (mm_interconnect_0_sd_card_avalon_sdcard_slave_read),                                    //                                                         .read
		.SD_Card_avalon_sdcard_slave_readdata                                (mm_interconnect_0_sd_card_avalon_sdcard_slave_readdata),                                //                                                         .readdata
		.SD_Card_avalon_sdcard_slave_writedata                               (mm_interconnect_0_sd_card_avalon_sdcard_slave_writedata),                               //                                                         .writedata
		.SD_Card_avalon_sdcard_slave_byteenable                              (mm_interconnect_0_sd_card_avalon_sdcard_slave_byteenable),                              //                                                         .byteenable
		.SD_Card_avalon_sdcard_slave_waitrequest                             (mm_interconnect_0_sd_card_avalon_sdcard_slave_waitrequest),                             //                                                         .waitrequest
		.SD_Card_avalon_sdcard_slave_chipselect                              (mm_interconnect_0_sd_card_avalon_sdcard_slave_chipselect),                              //                                                         .chipselect
		.SDRAM_s1_address                                                    (mm_interconnect_0_sdram_s1_address),                                                    //                                                 SDRAM_s1.address
		.SDRAM_s1_write                                                      (mm_interconnect_0_sdram_s1_write),                                                      //                                                         .write
		.SDRAM_s1_read                                                       (mm_interconnect_0_sdram_s1_read),                                                       //                                                         .read
		.SDRAM_s1_readdata                                                   (mm_interconnect_0_sdram_s1_readdata),                                                   //                                                         .readdata
		.SDRAM_s1_writedata                                                  (mm_interconnect_0_sdram_s1_writedata),                                                  //                                                         .writedata
		.SDRAM_s1_byteenable                                                 (mm_interconnect_0_sdram_s1_byteenable),                                                 //                                                         .byteenable
		.SDRAM_s1_readdatavalid                                              (mm_interconnect_0_sdram_s1_readdatavalid),                                              //                                                         .readdatavalid
		.SDRAM_s1_waitrequest                                                (mm_interconnect_0_sdram_s1_waitrequest),                                                //                                                         .waitrequest
		.SDRAM_s1_chipselect                                                 (mm_interconnect_0_sdram_s1_chipselect),                                                 //                                                         .chipselect
		.Serial_Port_avalon_rs232_slave_address                              (mm_interconnect_0_serial_port_avalon_rs232_slave_address),                              //                           Serial_Port_avalon_rs232_slave.address
		.Serial_Port_avalon_rs232_slave_write                                (mm_interconnect_0_serial_port_avalon_rs232_slave_write),                                //                                                         .write
		.Serial_Port_avalon_rs232_slave_read                                 (mm_interconnect_0_serial_port_avalon_rs232_slave_read),                                 //                                                         .read
		.Serial_Port_avalon_rs232_slave_readdata                             (mm_interconnect_0_serial_port_avalon_rs232_slave_readdata),                             //                                                         .readdata
		.Serial_Port_avalon_rs232_slave_writedata                            (mm_interconnect_0_serial_port_avalon_rs232_slave_writedata),                            //                                                         .writedata
		.Serial_Port_avalon_rs232_slave_byteenable                           (mm_interconnect_0_serial_port_avalon_rs232_slave_byteenable),                           //                                                         .byteenable
		.Serial_Port_avalon_rs232_slave_chipselect                           (mm_interconnect_0_serial_port_avalon_rs232_slave_chipselect),                           //                                                         .chipselect
		.Slider_Switches_s1_address                                          (mm_interconnect_0_slider_switches_s1_address),                                          //                                       Slider_Switches_s1.address
		.Slider_Switches_s1_readdata                                         (mm_interconnect_0_slider_switches_s1_readdata),                                         //                                                         .readdata
		.SRAM_avalon_sram_slave_address                                      (mm_interconnect_0_sram_avalon_sram_slave_address),                                      //                                   SRAM_avalon_sram_slave.address
		.SRAM_avalon_sram_slave_write                                        (mm_interconnect_0_sram_avalon_sram_slave_write),                                        //                                                         .write
		.SRAM_avalon_sram_slave_read                                         (mm_interconnect_0_sram_avalon_sram_slave_read),                                         //                                                         .read
		.SRAM_avalon_sram_slave_readdata                                     (mm_interconnect_0_sram_avalon_sram_slave_readdata),                                     //                                                         .readdata
		.SRAM_avalon_sram_slave_writedata                                    (mm_interconnect_0_sram_avalon_sram_slave_writedata),                                    //                                                         .writedata
		.SRAM_avalon_sram_slave_byteenable                                   (mm_interconnect_0_sram_avalon_sram_slave_byteenable),                                   //                                                         .byteenable
		.SRAM_avalon_sram_slave_readdatavalid                                (mm_interconnect_0_sram_avalon_sram_slave_readdatavalid),                                //                                                         .readdatavalid
		.SysID_control_slave_address                                         (mm_interconnect_0_sysid_control_slave_address),                                         //                                      SysID_control_slave.address
		.SysID_control_slave_readdata                                        (mm_interconnect_0_sysid_control_slave_readdata),                                        //                                                         .readdata
		.USB_avalon_usb_slave_address                                        (mm_interconnect_0_usb_avalon_usb_slave_address),                                        //                                     USB_avalon_usb_slave.address
		.USB_avalon_usb_slave_write                                          (mm_interconnect_0_usb_avalon_usb_slave_write),                                          //                                                         .write
		.USB_avalon_usb_slave_read                                           (mm_interconnect_0_usb_avalon_usb_slave_read),                                           //                                                         .read
		.USB_avalon_usb_slave_readdata                                       (mm_interconnect_0_usb_avalon_usb_slave_readdata),                                       //                                                         .readdata
		.USB_avalon_usb_slave_writedata                                      (mm_interconnect_0_usb_avalon_usb_slave_writedata),                                      //                                                         .writedata
		.USB_avalon_usb_slave_chipselect                                     (mm_interconnect_0_usb_avalon_usb_slave_chipselect),                                     //                                                         .chipselect
		.VGA_Subsystem_char_buffer_control_slave_address                     (mm_interconnect_0_vga_subsystem_char_buffer_control_slave_address),                     //                  VGA_Subsystem_char_buffer_control_slave.address
		.VGA_Subsystem_char_buffer_control_slave_write                       (mm_interconnect_0_vga_subsystem_char_buffer_control_slave_write),                       //                                                         .write
		.VGA_Subsystem_char_buffer_control_slave_read                        (mm_interconnect_0_vga_subsystem_char_buffer_control_slave_read),                        //                                                         .read
		.VGA_Subsystem_char_buffer_control_slave_readdata                    (mm_interconnect_0_vga_subsystem_char_buffer_control_slave_readdata),                    //                                                         .readdata
		.VGA_Subsystem_char_buffer_control_slave_writedata                   (mm_interconnect_0_vga_subsystem_char_buffer_control_slave_writedata),                   //                                                         .writedata
		.VGA_Subsystem_char_buffer_control_slave_byteenable                  (mm_interconnect_0_vga_subsystem_char_buffer_control_slave_byteenable),                  //                                                         .byteenable
		.VGA_Subsystem_char_buffer_slave_address                             (mm_interconnect_0_vga_subsystem_char_buffer_slave_address),                             //                          VGA_Subsystem_char_buffer_slave.address
		.VGA_Subsystem_char_buffer_slave_write                               (mm_interconnect_0_vga_subsystem_char_buffer_slave_write),                               //                                                         .write
		.VGA_Subsystem_char_buffer_slave_readdata                            (mm_interconnect_0_vga_subsystem_char_buffer_slave_readdata),                            //                                                         .readdata
		.VGA_Subsystem_char_buffer_slave_writedata                           (mm_interconnect_0_vga_subsystem_char_buffer_slave_writedata),                           //                                                         .writedata
		.VGA_Subsystem_char_buffer_slave_byteenable                          (mm_interconnect_0_vga_subsystem_char_buffer_slave_byteenable),                          //                                                         .byteenable
		.VGA_Subsystem_char_buffer_slave_chipselect                          (mm_interconnect_0_vga_subsystem_char_buffer_slave_chipselect),                          //                                                         .chipselect
		.VGA_Subsystem_char_buffer_slave_clken                               (mm_interconnect_0_vga_subsystem_char_buffer_slave_clken),                               //                                                         .clken
		.VGA_Subsystem_pixel_dma_control_slave_address                       (mm_interconnect_0_vga_subsystem_pixel_dma_control_slave_address),                       //                    VGA_Subsystem_pixel_dma_control_slave.address
		.VGA_Subsystem_pixel_dma_control_slave_write                         (mm_interconnect_0_vga_subsystem_pixel_dma_control_slave_write),                         //                                                         .write
		.VGA_Subsystem_pixel_dma_control_slave_read                          (mm_interconnect_0_vga_subsystem_pixel_dma_control_slave_read),                          //                                                         .read
		.VGA_Subsystem_pixel_dma_control_slave_readdata                      (mm_interconnect_0_vga_subsystem_pixel_dma_control_slave_readdata),                      //                                                         .readdata
		.VGA_Subsystem_pixel_dma_control_slave_writedata                     (mm_interconnect_0_vga_subsystem_pixel_dma_control_slave_writedata),                     //                                                         .writedata
		.VGA_Subsystem_pixel_dma_control_slave_byteenable                    (mm_interconnect_0_vga_subsystem_pixel_dma_control_slave_byteenable),                    //                                                         .byteenable
		.VGA_Subsystem_rgb_slave_read                                        (mm_interconnect_0_vga_subsystem_rgb_slave_read),                                        //                                  VGA_Subsystem_rgb_slave.read
		.VGA_Subsystem_rgb_slave_readdata                                    (mm_interconnect_0_vga_subsystem_rgb_slave_readdata),                                    //                                                         .readdata
		.Video_In_Subsystem_video_in_dma_control_slave_address               (mm_interconnect_0_video_in_subsystem_video_in_dma_control_slave_address),               //            Video_In_Subsystem_video_in_dma_control_slave.address
		.Video_In_Subsystem_video_in_dma_control_slave_write                 (mm_interconnect_0_video_in_subsystem_video_in_dma_control_slave_write),                 //                                                         .write
		.Video_In_Subsystem_video_in_dma_control_slave_read                  (mm_interconnect_0_video_in_subsystem_video_in_dma_control_slave_read),                  //                                                         .read
		.Video_In_Subsystem_video_in_dma_control_slave_readdata              (mm_interconnect_0_video_in_subsystem_video_in_dma_control_slave_readdata),              //                                                         .readdata
		.Video_In_Subsystem_video_in_dma_control_slave_writedata             (mm_interconnect_0_video_in_subsystem_video_in_dma_control_slave_writedata),             //                                                         .writedata
		.Video_In_Subsystem_video_in_dma_control_slave_byteenable            (mm_interconnect_0_video_in_subsystem_video_in_dma_control_slave_byteenable),            //                                                         .byteenable
		.Video_In_Subsystem_video_in_edge_detection_control_slave_address    (mm_interconnect_0_video_in_subsystem_video_in_edge_detection_control_slave_address),    // Video_In_Subsystem_video_in_edge_detection_control_slave.address
		.Video_In_Subsystem_video_in_edge_detection_control_slave_write      (mm_interconnect_0_video_in_subsystem_video_in_edge_detection_control_slave_write),      //                                                         .write
		.Video_In_Subsystem_video_in_edge_detection_control_slave_readdata   (mm_interconnect_0_video_in_subsystem_video_in_edge_detection_control_slave_readdata),   //                                                         .readdata
		.Video_In_Subsystem_video_in_edge_detection_control_slave_writedata  (mm_interconnect_0_video_in_subsystem_video_in_edge_detection_control_slave_writedata),  //                                                         .writedata
		.Video_In_Subsystem_video_in_edge_detection_control_slave_chipselect (mm_interconnect_0_video_in_subsystem_video_in_edge_detection_control_slave_chipselect)  //                                                         .chipselect
	);

	Computer_System_irq_mapper irq_mapper (
		.clk            (system_pll_sys_clk_clk),             //        clk.clk
		.reset          (rst_controller_001_reset_out_reset), //  clk_reset.reset
		.receiver0_irq  (irq_mapper_receiver0_irq),           //  receiver0.irq
		.receiver1_irq  (irq_mapper_receiver1_irq),           //  receiver1.irq
		.receiver2_irq  (irq_mapper_receiver2_irq),           //  receiver2.irq
		.receiver3_irq  (irq_mapper_receiver3_irq),           //  receiver3.irq
		.receiver4_irq  (irq_mapper_receiver4_irq),           //  receiver4.irq
		.receiver5_irq  (irq_mapper_receiver5_irq),           //  receiver5.irq
		.receiver6_irq  (irq_mapper_receiver6_irq),           //  receiver6.irq
		.receiver7_irq  (irq_mapper_receiver7_irq),           //  receiver7.irq
		.receiver8_irq  (irq_mapper_receiver8_irq),           //  receiver8.irq
		.receiver9_irq  (irq_mapper_receiver9_irq),           //  receiver9.irq
		.receiver10_irq (irq_mapper_receiver10_irq),          // receiver10.irq
		.sender_irq     (nios2_irq_irq)                       //     sender.irq
	);

	Computer_System_irq_mapper irq_mapper_001 (
		.clk            (system_pll_sys_clk_clk),             //        clk.clk
		.reset          (rst_controller_002_reset_out_reset), //  clk_reset.reset
		.receiver0_irq  (irq_mapper_receiver0_irq),           //  receiver0.irq
		.receiver1_irq  (irq_mapper_receiver1_irq),           //  receiver1.irq
		.receiver2_irq  (irq_mapper_receiver2_irq),           //  receiver2.irq
		.receiver3_irq  (irq_mapper_receiver3_irq),           //  receiver3.irq
		.receiver4_irq  (irq_mapper_receiver4_irq),           //  receiver4.irq
		.receiver5_irq  (irq_mapper_receiver5_irq),           //  receiver5.irq
		.receiver6_irq  (irq_mapper_receiver6_irq),           //  receiver6.irq
		.receiver7_irq  (irq_mapper_receiver7_irq),           //  receiver7.irq
		.receiver8_irq  (irq_mapper_001_receiver8_irq),       //  receiver8.irq
		.receiver9_irq  (irq_mapper_001_receiver9_irq),       //  receiver9.irq
		.receiver10_irq (irq_mapper_001_receiver10_irq),      // receiver10.irq
		.sender_irq     (nios2_2nd_core_irq_irq)              //     sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (system_pll_reset_source_reset),  // reset_in0.reset
		.clk            (system_pll_sys_clk_clk),         //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (nios2_debug_reset_request_reset),    // reset_in0.reset
		.reset_in1      (system_pll_reset_source_reset),      // reset_in1.reset
		.clk            (system_pll_sys_clk_clk),             //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (nios2_2nd_core_debug_reset_request_reset), // reset_in0.reset
		.reset_in1      (system_pll_reset_source_reset),            // reset_in1.reset
		.clk            (system_pll_sys_clk_clk),                   //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset),       // reset_out.reset
		.reset_req      (),                                         // (terminated)
		.reset_req_in0  (1'b0),                                     // (terminated)
		.reset_req_in1  (1'b0),                                     // (terminated)
		.reset_in2      (1'b0),                                     // (terminated)
		.reset_req_in2  (1'b0),                                     // (terminated)
		.reset_in3      (1'b0),                                     // (terminated)
		.reset_req_in3  (1'b0),                                     // (terminated)
		.reset_in4      (1'b0),                                     // (terminated)
		.reset_req_in4  (1'b0),                                     // (terminated)
		.reset_in5      (1'b0),                                     // (terminated)
		.reset_req_in5  (1'b0),                                     // (terminated)
		.reset_in6      (1'b0),                                     // (terminated)
		.reset_req_in6  (1'b0),                                     // (terminated)
		.reset_in7      (1'b0),                                     // (terminated)
		.reset_req_in7  (1'b0),                                     // (terminated)
		.reset_in8      (1'b0),                                     // (terminated)
		.reset_req_in8  (1'b0),                                     // (terminated)
		.reset_in9      (1'b0),                                     // (terminated)
		.reset_req_in9  (1'b0),                                     // (terminated)
		.reset_in10     (1'b0),                                     // (terminated)
		.reset_req_in10 (1'b0),                                     // (terminated)
		.reset_in11     (1'b0),                                     // (terminated)
		.reset_req_in11 (1'b0),                                     // (terminated)
		.reset_in12     (1'b0),                                     // (terminated)
		.reset_req_in12 (1'b0),                                     // (terminated)
		.reset_in13     (1'b0),                                     // (terminated)
		.reset_req_in13 (1'b0),                                     // (terminated)
		.reset_in14     (1'b0),                                     // (terminated)
		.reset_req_in14 (1'b0),                                     // (terminated)
		.reset_in15     (1'b0),                                     // (terminated)
		.reset_req_in15 (1'b0)                                      // (terminated)
	);

endmodule
